VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aes_core
  CLASS BLOCK ;
  FOREIGN aes_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1242.000 BY 1259.920 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 1255.920 733.040 1258.920 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 1255.920 161.840 1258.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 947.520 4.000 948.080 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1246.560 1241.000 1247.120 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 1255.920 914.480 1258.920 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 809.760 1241.000 810.320 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 581.280 4.000 581.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 456.960 1241.000 457.520 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1249.920 4.000 1250.480 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1216.320 1255.920 1216.880 1258.920 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 994.560 4.000 995.120 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 201.600 1241.000 202.160 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 641.760 4.000 642.320 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1255.920 269.360 1258.920 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1115.520 4.000 1116.080 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 1.000 1069.040 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 262.080 1241.000 262.640 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1212.960 1.000 1213.520 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.480 4.000 61.040 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1229.760 1255.920 1230.320 1258.920 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1255.920 635.600 1258.920 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 131.040 4.000 131.600 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 241.920 4.000 242.480 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1255.920 598.640 1258.920 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1209.600 1241.000 1210.160 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1255.920 134.960 1258.920 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 940.800 1241.000 941.360 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 715.680 4.000 716.240 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 1255.920 1058.960 1258.920 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 309.120 1241.000 309.680 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 436.800 4.000 437.360 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 530.880 1241.000 531.440 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 1255.920 101.360 1258.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1011.360 1255.920 1011.920 1258.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1.000 437.360 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 967.680 1241.000 968.240 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 1.000 252.560 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 117.600 1241.000 118.160 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 211.680 1241.000 212.240 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 1.000 921.200 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 1255.920 682.640 1258.920 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1212.960 4.000 1213.520 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 23.520 4.000 24.080 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 1255.920 208.880 1258.920 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1255.920 329.840 1258.920 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1255.920 171.920 1258.920 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 934.080 4.000 934.640 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 1.000 739.760 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1088.640 1241.000 1089.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 275.520 1241.000 276.080 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 957.600 4.000 958.160 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 1.000 1166.480 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1078.560 4.000 1079.120 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 1.000 1032.080 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1255.920 538.160 1258.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 1255.920 672.560 1258.920 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1115.520 1.000 1116.080 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 443.520 1241.000 444.080 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 900.480 1255.920 901.040 1258.920 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1048.320 1255.920 1048.880 1258.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 1.000 121.520 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1179.360 1255.920 1179.920 1258.920 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 1.000 497.840 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 1255.920 185.360 1258.920 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 1255.920 50.960 1258.920 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 557.760 4.000 558.320 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 1.000 1045.520 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 493.920 1241.000 494.480 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 1255.920 1095.920 1258.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 423.360 4.000 423.920 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 188.160 1241.000 188.720 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1145.760 1255.920 1146.320 1258.920 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1.000 521.360 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1.000 776.720 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 141.120 1241.000 141.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 782.880 1241.000 783.440 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 850.080 4.000 850.640 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1135.680 1241.000 1136.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 1255.920 561.680 1258.920 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1.000 145.040 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 836.640 4.000 837.200 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 1.000 800.240 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 712.320 1241.000 712.880 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 1.000 558.320 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 1.000 410.480 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 406.560 1241.000 407.120 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 1.000 1055.600 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 507.360 4.000 507.920 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1169.280 1255.920 1169.840 1258.920 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1236.480 4.000 1237.040 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 655.200 4.000 655.760 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 1.000 823.760 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 1255.920 706.160 1258.920 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 789.600 4.000 790.160 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 248.640 1241.000 249.200 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.760 4.000 474.320 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 567.840 4.000 568.400 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 1.000 813.680 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 178.080 1241.000 178.640 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1233.120 1241.000 1233.680 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 43.680 1241.000 44.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1255.920 282.800 1258.920 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1255.920 608.720 1258.920 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 520.800 4.000 521.360 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 725.760 4.000 726.320 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 766.080 1255.920 766.640 1258.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 1.000 897.680 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 1255.920 111.440 1258.920 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 376.320 4.000 376.880 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1226.400 1.000 1226.960 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 1.000 460.880 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 1.000 376.880 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 1255.920 514.640 1258.920 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 1255.920 1132.880 1258.920 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 1.000 581.840 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 762.720 4.000 763.280 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 1255.920 974.960 1258.920 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1223.040 1241.000 1223.600 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 322.560 1241.000 323.120 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 813.120 4.000 813.680 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 238.560 1241.000 239.120 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.960 4.000 121.520 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.560 4.000 71.120 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 1255.920 998.480 1258.920 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 1255.920 780.080 1258.920 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1038.240 1241.000 1038.800 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 1255.920 924.560 1258.920 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 604.800 4.000 605.360 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1068.480 4.000 1069.040 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1149.120 1241.000 1149.680 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 688.800 1241.000 689.360 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1226.400 4.000 1226.960 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 517.440 1241.000 518.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1075.200 1241.000 1075.760 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1176.000 1.000 1176.560 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.960 4.000 289.520 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 873.600 1.000 874.160 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 1255.920 450.800 1258.920 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 860.160 4.000 860.720 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 1255.920 524.720 1258.920 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 1255.920 840.560 1258.920 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 1.000 423.920 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 1.000 595.280 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1189.440 4.000 1190.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 534.240 4.000 534.800 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 887.040 4.000 887.600 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 907.200 1241.000 907.760 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 893.760 1241.000 894.320 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.520 4.000 108.080 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 325.920 4.000 326.480 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 94.080 4.000 94.640 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1255.920 501.200 1258.920 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 1.000 568.400 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1139.040 4.000 1139.600 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 1255.920 380.240 1258.920 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 336.000 1241.000 336.560 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 339.360 4.000 339.920 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 349.440 4.000 350.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 30.240 1241.000 30.800 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 1.000 447.440 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 483.840 4.000 484.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 1.000 218.960 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 1255.920 864.080 1258.920 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 1255.920 951.440 1258.920 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 1.000 726.320 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 601.440 1241.000 602.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 618.240 4.000 618.800 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 1255.920 3.920 1258.920 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1044.960 4.000 1045.520 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 1255.920 696.080 1258.920 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.440 4.000 182.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 776.160 4.000 776.720 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 1.000 887.600 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 910.560 4.000 911.120 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 1255.920 353.360 1258.920 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 504.000 1241.000 504.560 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1172.640 1241.000 1173.200 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 675.360 1241.000 675.920 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1255.920 622.160 1258.920 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 1255.920 548.240 1258.920 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 1.000 655.760 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 577.920 1241.000 578.480 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 1255.920 585.200 1258.920 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 870.240 1241.000 870.800 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 1255.920 659.120 1258.920 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.520 4.000 192.080 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 1255.920 1082.480 1258.920 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1.000 168.560 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 168.000 4.000 168.560 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 1.000 534.800 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 981.120 4.000 981.680 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 564.480 1241.000 565.040 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 1255.920 37.520 1258.920 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1255.920 195.440 1258.920 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1255.920 27.440 1258.920 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 1.000 605.360 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 1.000 339.920 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1004.640 1241.000 1005.200 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 480.480 1241.000 481.040 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 20.160 1241.000 20.720 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 164.640 1241.000 165.200 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 1255.920 877.520 1258.920 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1128.960 4.000 1129.520 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 369.600 1241.000 370.160 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1051.680 1241.000 1052.240 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1.000 71.120 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 1.000 507.920 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 1255.920 756.560 1258.920 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 1.000 1139.600 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 897.120 4.000 897.680 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1.000 289.520 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 1.000 1129.520 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 1255.920 719.600 1258.920 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 1255.920 440.720 1258.920 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 460.320 4.000 460.880 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 80.640 1241.000 81.200 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1.000 692.720 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1176.000 4.000 1176.560 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 1255.920 477.680 1258.920 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 285.600 1241.000 286.160 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1008.000 4.000 1008.560 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 856.800 1241.000 857.360 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1112.160 1241.000 1112.720 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 749.280 1241.000 749.840 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1021.440 1255.920 1022.000 1258.920 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 1.000 326.480 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1078.560 1.000 1079.120 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 90.720 1241.000 91.280 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 873.600 4.000 874.160 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1206.240 1255.920 1206.800 1258.920 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1165.920 4.000 1166.480 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 591.360 1241.000 591.920 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 467.040 1241.000 467.600 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 880.320 1241.000 880.880 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 698.880 1241.000 699.440 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 1255.920 487.760 1258.920 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 446.880 4.000 447.440 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 47.040 4.000 47.600 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 1.000 1092.560 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1.000 182.000 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 157.920 4.000 158.480 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 1255.920 87.920 1258.920 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 104.160 1241.000 104.720 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 1255.920 245.840 1258.920 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1105.440 4.000 1106.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1255.920 222.320 1258.920 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.600 4.000 34.160 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1.000 350.000 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.840 4.000 316.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1105.440 1.000 1106.000 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1255.920 259.280 1258.920 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 651.840 1241.000 652.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1186.080 1241.000 1186.640 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1239.840 1255.920 1240.400 1258.920 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1065.120 1241.000 1065.680 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1028.160 1241.000 1028.720 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1014.720 1241.000 1015.280 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 1.000 632.240 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 1255.920 1119.440 1258.920 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1.000 34.160 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 1.000 10.640 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 1255.920 14.000 1258.920 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 1.000 642.320 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.320 4.000 544.880 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 692.160 4.000 692.720 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1255.920 464.240 1258.920 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 799.680 4.000 800.240 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 1.000 242.480 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1.000 544.880 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 631.680 4.000 632.240 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 1.000 995.120 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1.000 474.320 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 920.640 4.000 921.200 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 614.880 1241.000 615.440 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 833.280 1241.000 833.840 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 1.000 958.160 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 1255.920 403.760 1258.920 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1236.480 1.000 1237.040 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 796.320 1241.000 796.880 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 752.640 4.000 753.200 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 638.400 1241.000 638.960 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 1.000 948.080 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1108.800 1255.920 1109.360 1258.920 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 127.680 1241.000 128.240 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 1255.920 743.120 1258.920 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 1.000 1153.040 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 1255.920 306.320 1258.920 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1.000 158.480 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 10.080 4.000 10.640 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1202.880 4.000 1203.440 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 819.840 1241.000 820.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1.000 316.400 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1189.440 1.000 1190.000 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 1255.920 1072.400 1258.920 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 954.240 1241.000 954.800 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 1255.920 319.760 1258.920 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1255.920 427.280 1258.920 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1242.940 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1242.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1242.940 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 225.120 1241.000 225.680 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 1255.920 232.400 1258.920 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 433.440 1241.000 434.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 1255.920 830.480 1258.920 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 1255.920 575.120 1258.920 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 1255.920 74.480 1258.920 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1.000 108.080 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 917.280 1241.000 917.840 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 846.720 1241.000 847.280 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1.000 790.160 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 702.240 4.000 702.800 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 396.480 1241.000 397.040 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1202.880 1.000 1203.440 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 1255.920 803.600 1258.920 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 1.000 702.800 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1008.000 1.000 1008.560 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 299.040 1241.000 299.600 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 1255.920 148.400 1258.920 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.400 4.000 218.960 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 1.000 131.600 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 1255.920 417.200 1258.920 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 735.840 1241.000 736.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1196.160 1241.000 1196.720 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.480 4.000 145.040 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 497.280 4.000 497.840 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 540.960 1241.000 541.520 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 1.000 971.600 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 1255.920 961.520 1258.920 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 1.000 934.640 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 1.000 61.040 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 6.720 1241.000 7.280 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 346.080 1241.000 346.640 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 1255.920 390.320 1258.920 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1098.720 1241.000 1099.280 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 971.040 4.000 971.600 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1055.040 4.000 1055.600 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1018.080 4.000 1018.640 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 1.000 47.600 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 265.440 4.000 266.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 661.920 1241.000 662.480 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 1.000 716.240 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.960 4.000 205.520 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1155.840 1255.920 1156.400 1258.920 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 1255.920 64.400 1258.920 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1.000 192.080 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 759.360 1241.000 759.920 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 1255.920 1193.360 1258.920 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 739.200 4.000 739.760 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 991.200 1241.000 991.760 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 420.000 1241.000 420.560 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 1.000 860.720 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1034.880 1255.920 1035.440 1258.920 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 1255.920 292.880 1258.920 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1.000 386.960 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 772.800 1241.000 773.360 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 1.000 1018.640 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 383.040 1241.000 383.600 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 53.760 1241.000 54.320 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1.000 205.520 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 1.000 618.800 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 554.400 1241.000 554.960 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 987.840 1255.920 988.400 1258.920 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1125.600 1241.000 1126.160 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 67.200 1241.000 67.760 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 252.000 4.000 252.560 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 722.400 1241.000 722.960 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1.000 24.080 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 1162.560 1241.000 1163.120 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 1255.920 938.000 1258.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 151.200 1241.000 151.760 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 1255.920 890.960 1258.920 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 1.000 850.640 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.400 4.000 386.960 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 1.000 837.200 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 1.000 981.680 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 594.720 4.000 595.280 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1092.000 4.000 1092.560 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 1255.920 343.280 1258.920 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 409.920 4.000 410.480 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 1.000 266.000 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1.000 94.640 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1255.920 645.680 1258.920 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 1255.920 366.800 1258.920 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1.000 679.280 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 1255.920 854.000 1258.920 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 359.520 1241.000 360.080 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 823.200 4.000 823.760 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 977.760 1241.000 978.320 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 1.000 279.440 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1.000 484.400 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 1.000 753.200 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 930.720 1241.000 931.280 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 1.000 763.280 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 1255.920 817.040 1258.920 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 1255.920 793.520 1258.920 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1152.480 4.000 1153.040 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1255.920 124.880 1258.920 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 1.000 911.120 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 278.880 4.000 279.440 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1031.520 4.000 1032.080 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1238.000 624.960 1241.000 625.520 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 1234.800 1242.940 ;
      LAYER Metal2 ;
        RECT 0.140 1255.620 3.060 1256.500 ;
        RECT 4.220 1255.620 13.140 1256.500 ;
        RECT 14.300 1255.620 26.580 1256.500 ;
        RECT 27.740 1255.620 36.660 1256.500 ;
        RECT 37.820 1255.620 50.100 1256.500 ;
        RECT 51.260 1255.620 63.540 1256.500 ;
        RECT 64.700 1255.620 73.620 1256.500 ;
        RECT 74.780 1255.620 87.060 1256.500 ;
        RECT 88.220 1255.620 100.500 1256.500 ;
        RECT 101.660 1255.620 110.580 1256.500 ;
        RECT 111.740 1255.620 124.020 1256.500 ;
        RECT 125.180 1255.620 134.100 1256.500 ;
        RECT 135.260 1255.620 147.540 1256.500 ;
        RECT 148.700 1255.620 160.980 1256.500 ;
        RECT 162.140 1255.620 171.060 1256.500 ;
        RECT 172.220 1255.620 184.500 1256.500 ;
        RECT 185.660 1255.620 194.580 1256.500 ;
        RECT 195.740 1255.620 208.020 1256.500 ;
        RECT 209.180 1255.620 221.460 1256.500 ;
        RECT 222.620 1255.620 231.540 1256.500 ;
        RECT 232.700 1255.620 244.980 1256.500 ;
        RECT 246.140 1255.620 258.420 1256.500 ;
        RECT 259.580 1255.620 268.500 1256.500 ;
        RECT 269.660 1255.620 281.940 1256.500 ;
        RECT 283.100 1255.620 292.020 1256.500 ;
        RECT 293.180 1255.620 305.460 1256.500 ;
        RECT 306.620 1255.620 318.900 1256.500 ;
        RECT 320.060 1255.620 328.980 1256.500 ;
        RECT 330.140 1255.620 342.420 1256.500 ;
        RECT 343.580 1255.620 352.500 1256.500 ;
        RECT 353.660 1255.620 365.940 1256.500 ;
        RECT 367.100 1255.620 379.380 1256.500 ;
        RECT 380.540 1255.620 389.460 1256.500 ;
        RECT 390.620 1255.620 402.900 1256.500 ;
        RECT 404.060 1255.620 416.340 1256.500 ;
        RECT 417.500 1255.620 426.420 1256.500 ;
        RECT 427.580 1255.620 439.860 1256.500 ;
        RECT 441.020 1255.620 449.940 1256.500 ;
        RECT 451.100 1255.620 463.380 1256.500 ;
        RECT 464.540 1255.620 476.820 1256.500 ;
        RECT 477.980 1255.620 486.900 1256.500 ;
        RECT 488.060 1255.620 500.340 1256.500 ;
        RECT 501.500 1255.620 513.780 1256.500 ;
        RECT 514.940 1255.620 523.860 1256.500 ;
        RECT 525.020 1255.620 537.300 1256.500 ;
        RECT 538.460 1255.620 547.380 1256.500 ;
        RECT 548.540 1255.620 560.820 1256.500 ;
        RECT 561.980 1255.620 574.260 1256.500 ;
        RECT 575.420 1255.620 584.340 1256.500 ;
        RECT 585.500 1255.620 597.780 1256.500 ;
        RECT 598.940 1255.620 607.860 1256.500 ;
        RECT 609.020 1255.620 621.300 1256.500 ;
        RECT 622.460 1255.620 634.740 1256.500 ;
        RECT 635.900 1255.620 644.820 1256.500 ;
        RECT 645.980 1255.620 658.260 1256.500 ;
        RECT 659.420 1255.620 671.700 1256.500 ;
        RECT 672.860 1255.620 681.780 1256.500 ;
        RECT 682.940 1255.620 695.220 1256.500 ;
        RECT 696.380 1255.620 705.300 1256.500 ;
        RECT 706.460 1255.620 718.740 1256.500 ;
        RECT 719.900 1255.620 732.180 1256.500 ;
        RECT 733.340 1255.620 742.260 1256.500 ;
        RECT 743.420 1255.620 755.700 1256.500 ;
        RECT 756.860 1255.620 765.780 1256.500 ;
        RECT 766.940 1255.620 779.220 1256.500 ;
        RECT 780.380 1255.620 792.660 1256.500 ;
        RECT 793.820 1255.620 802.740 1256.500 ;
        RECT 803.900 1255.620 816.180 1256.500 ;
        RECT 817.340 1255.620 829.620 1256.500 ;
        RECT 830.780 1255.620 839.700 1256.500 ;
        RECT 840.860 1255.620 853.140 1256.500 ;
        RECT 854.300 1255.620 863.220 1256.500 ;
        RECT 864.380 1255.620 876.660 1256.500 ;
        RECT 877.820 1255.620 890.100 1256.500 ;
        RECT 891.260 1255.620 900.180 1256.500 ;
        RECT 901.340 1255.620 913.620 1256.500 ;
        RECT 914.780 1255.620 923.700 1256.500 ;
        RECT 924.860 1255.620 937.140 1256.500 ;
        RECT 938.300 1255.620 950.580 1256.500 ;
        RECT 951.740 1255.620 960.660 1256.500 ;
        RECT 961.820 1255.620 974.100 1256.500 ;
        RECT 975.260 1255.620 987.540 1256.500 ;
        RECT 988.700 1255.620 997.620 1256.500 ;
        RECT 998.780 1255.620 1011.060 1256.500 ;
        RECT 1012.220 1255.620 1021.140 1256.500 ;
        RECT 1022.300 1255.620 1034.580 1256.500 ;
        RECT 1035.740 1255.620 1048.020 1256.500 ;
        RECT 1049.180 1255.620 1058.100 1256.500 ;
        RECT 1059.260 1255.620 1071.540 1256.500 ;
        RECT 1072.700 1255.620 1081.620 1256.500 ;
        RECT 1082.780 1255.620 1095.060 1256.500 ;
        RECT 1096.220 1255.620 1108.500 1256.500 ;
        RECT 1109.660 1255.620 1118.580 1256.500 ;
        RECT 1119.740 1255.620 1132.020 1256.500 ;
        RECT 1133.180 1255.620 1145.460 1256.500 ;
        RECT 1146.620 1255.620 1155.540 1256.500 ;
        RECT 1156.700 1255.620 1168.980 1256.500 ;
        RECT 1170.140 1255.620 1179.060 1256.500 ;
        RECT 1180.220 1255.620 1192.500 1256.500 ;
        RECT 1193.660 1255.620 1205.940 1256.500 ;
        RECT 1207.100 1255.620 1216.020 1256.500 ;
        RECT 1217.180 1255.620 1229.460 1256.500 ;
        RECT 1230.620 1255.620 1235.780 1256.500 ;
        RECT 0.140 4.300 1235.780 1255.620 ;
        RECT 0.860 4.000 9.780 4.300 ;
        RECT 10.940 4.000 23.220 4.300 ;
        RECT 24.380 4.000 33.300 4.300 ;
        RECT 34.460 4.000 46.740 4.300 ;
        RECT 47.900 4.000 60.180 4.300 ;
        RECT 61.340 4.000 70.260 4.300 ;
        RECT 71.420 4.000 83.700 4.300 ;
        RECT 84.860 4.000 93.780 4.300 ;
        RECT 94.940 4.000 107.220 4.300 ;
        RECT 108.380 4.000 120.660 4.300 ;
        RECT 121.820 4.000 130.740 4.300 ;
        RECT 131.900 4.000 144.180 4.300 ;
        RECT 145.340 4.000 157.620 4.300 ;
        RECT 158.780 4.000 167.700 4.300 ;
        RECT 168.860 4.000 181.140 4.300 ;
        RECT 182.300 4.000 191.220 4.300 ;
        RECT 192.380 4.000 204.660 4.300 ;
        RECT 205.820 4.000 218.100 4.300 ;
        RECT 219.260 4.000 228.180 4.300 ;
        RECT 229.340 4.000 241.620 4.300 ;
        RECT 242.780 4.000 251.700 4.300 ;
        RECT 252.860 4.000 265.140 4.300 ;
        RECT 266.300 4.000 278.580 4.300 ;
        RECT 279.740 4.000 288.660 4.300 ;
        RECT 289.820 4.000 302.100 4.300 ;
        RECT 303.260 4.000 315.540 4.300 ;
        RECT 316.700 4.000 325.620 4.300 ;
        RECT 326.780 4.000 339.060 4.300 ;
        RECT 340.220 4.000 349.140 4.300 ;
        RECT 350.300 4.000 362.580 4.300 ;
        RECT 363.740 4.000 376.020 4.300 ;
        RECT 377.180 4.000 386.100 4.300 ;
        RECT 387.260 4.000 399.540 4.300 ;
        RECT 400.700 4.000 409.620 4.300 ;
        RECT 410.780 4.000 423.060 4.300 ;
        RECT 424.220 4.000 436.500 4.300 ;
        RECT 437.660 4.000 446.580 4.300 ;
        RECT 447.740 4.000 460.020 4.300 ;
        RECT 461.180 4.000 473.460 4.300 ;
        RECT 474.620 4.000 483.540 4.300 ;
        RECT 484.700 4.000 496.980 4.300 ;
        RECT 498.140 4.000 507.060 4.300 ;
        RECT 508.220 4.000 520.500 4.300 ;
        RECT 521.660 4.000 533.940 4.300 ;
        RECT 535.100 4.000 544.020 4.300 ;
        RECT 545.180 4.000 557.460 4.300 ;
        RECT 558.620 4.000 567.540 4.300 ;
        RECT 568.700 4.000 580.980 4.300 ;
        RECT 582.140 4.000 594.420 4.300 ;
        RECT 595.580 4.000 604.500 4.300 ;
        RECT 605.660 4.000 617.940 4.300 ;
        RECT 619.100 4.000 631.380 4.300 ;
        RECT 632.540 4.000 641.460 4.300 ;
        RECT 642.620 4.000 654.900 4.300 ;
        RECT 656.060 4.000 664.980 4.300 ;
        RECT 666.140 4.000 678.420 4.300 ;
        RECT 679.580 4.000 691.860 4.300 ;
        RECT 693.020 4.000 701.940 4.300 ;
        RECT 703.100 4.000 715.380 4.300 ;
        RECT 716.540 4.000 725.460 4.300 ;
        RECT 726.620 4.000 738.900 4.300 ;
        RECT 740.060 4.000 752.340 4.300 ;
        RECT 753.500 4.000 762.420 4.300 ;
        RECT 763.580 4.000 775.860 4.300 ;
        RECT 777.020 4.000 789.300 4.300 ;
        RECT 790.460 4.000 799.380 4.300 ;
        RECT 800.540 4.000 812.820 4.300 ;
        RECT 813.980 4.000 822.900 4.300 ;
        RECT 824.060 4.000 836.340 4.300 ;
        RECT 837.500 4.000 849.780 4.300 ;
        RECT 850.940 4.000 859.860 4.300 ;
        RECT 861.020 4.000 873.300 4.300 ;
        RECT 874.460 4.000 886.740 4.300 ;
        RECT 887.900 4.000 896.820 4.300 ;
        RECT 897.980 4.000 910.260 4.300 ;
        RECT 911.420 4.000 920.340 4.300 ;
        RECT 921.500 4.000 933.780 4.300 ;
        RECT 934.940 4.000 947.220 4.300 ;
        RECT 948.380 4.000 957.300 4.300 ;
        RECT 958.460 4.000 970.740 4.300 ;
        RECT 971.900 4.000 980.820 4.300 ;
        RECT 981.980 4.000 994.260 4.300 ;
        RECT 995.420 4.000 1007.700 4.300 ;
        RECT 1008.860 4.000 1017.780 4.300 ;
        RECT 1018.940 4.000 1031.220 4.300 ;
        RECT 1032.380 4.000 1044.660 4.300 ;
        RECT 1045.820 4.000 1054.740 4.300 ;
        RECT 1055.900 4.000 1068.180 4.300 ;
        RECT 1069.340 4.000 1078.260 4.300 ;
        RECT 1079.420 4.000 1091.700 4.300 ;
        RECT 1092.860 4.000 1105.140 4.300 ;
        RECT 1106.300 4.000 1115.220 4.300 ;
        RECT 1116.380 4.000 1128.660 4.300 ;
        RECT 1129.820 4.000 1138.740 4.300 ;
        RECT 1139.900 4.000 1152.180 4.300 ;
        RECT 1153.340 4.000 1165.620 4.300 ;
        RECT 1166.780 4.000 1175.700 4.300 ;
        RECT 1176.860 4.000 1189.140 4.300 ;
        RECT 1190.300 4.000 1202.580 4.300 ;
        RECT 1203.740 4.000 1212.660 4.300 ;
        RECT 1213.820 4.000 1226.100 4.300 ;
        RECT 1227.260 4.000 1235.780 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 1237.340 1241.940 1244.740 ;
        RECT 0.090 1236.180 0.700 1237.340 ;
        RECT 4.300 1236.180 1241.940 1237.340 ;
        RECT 0.090 1233.980 1241.940 1236.180 ;
        RECT 0.090 1232.820 1237.700 1233.980 ;
        RECT 1241.300 1232.820 1241.940 1233.980 ;
        RECT 0.090 1227.260 1241.940 1232.820 ;
        RECT 0.090 1226.100 0.700 1227.260 ;
        RECT 4.300 1226.100 1241.940 1227.260 ;
        RECT 0.090 1223.900 1241.940 1226.100 ;
        RECT 0.090 1222.740 1237.700 1223.900 ;
        RECT 1241.300 1222.740 1241.940 1223.900 ;
        RECT 0.090 1213.820 1241.940 1222.740 ;
        RECT 0.090 1212.660 0.700 1213.820 ;
        RECT 4.300 1212.660 1241.940 1213.820 ;
        RECT 0.090 1210.460 1241.940 1212.660 ;
        RECT 0.090 1209.300 1237.700 1210.460 ;
        RECT 1241.300 1209.300 1241.940 1210.460 ;
        RECT 0.090 1203.740 1241.940 1209.300 ;
        RECT 0.090 1202.580 0.700 1203.740 ;
        RECT 4.300 1202.580 1241.940 1203.740 ;
        RECT 0.090 1197.020 1241.940 1202.580 ;
        RECT 0.090 1195.860 1237.700 1197.020 ;
        RECT 1241.300 1195.860 1241.940 1197.020 ;
        RECT 0.090 1190.300 1241.940 1195.860 ;
        RECT 0.090 1189.140 0.700 1190.300 ;
        RECT 4.300 1189.140 1241.940 1190.300 ;
        RECT 0.090 1186.940 1241.940 1189.140 ;
        RECT 0.090 1185.780 1237.700 1186.940 ;
        RECT 1241.300 1185.780 1241.940 1186.940 ;
        RECT 0.090 1176.860 1241.940 1185.780 ;
        RECT 0.090 1175.700 0.700 1176.860 ;
        RECT 4.300 1175.700 1241.940 1176.860 ;
        RECT 0.090 1173.500 1241.940 1175.700 ;
        RECT 0.090 1172.340 1237.700 1173.500 ;
        RECT 1241.300 1172.340 1241.940 1173.500 ;
        RECT 0.090 1166.780 1241.940 1172.340 ;
        RECT 0.090 1165.620 0.700 1166.780 ;
        RECT 4.300 1165.620 1241.940 1166.780 ;
        RECT 0.090 1163.420 1241.940 1165.620 ;
        RECT 0.090 1162.260 1237.700 1163.420 ;
        RECT 1241.300 1162.260 1241.940 1163.420 ;
        RECT 0.090 1153.340 1241.940 1162.260 ;
        RECT 0.090 1152.180 0.700 1153.340 ;
        RECT 4.300 1152.180 1241.940 1153.340 ;
        RECT 0.090 1149.980 1241.940 1152.180 ;
        RECT 0.090 1148.820 1237.700 1149.980 ;
        RECT 1241.300 1148.820 1241.940 1149.980 ;
        RECT 0.090 1139.900 1241.940 1148.820 ;
        RECT 0.090 1138.740 0.700 1139.900 ;
        RECT 4.300 1138.740 1241.940 1139.900 ;
        RECT 0.090 1136.540 1241.940 1138.740 ;
        RECT 0.090 1135.380 1237.700 1136.540 ;
        RECT 1241.300 1135.380 1241.940 1136.540 ;
        RECT 0.090 1129.820 1241.940 1135.380 ;
        RECT 0.090 1128.660 0.700 1129.820 ;
        RECT 4.300 1128.660 1241.940 1129.820 ;
        RECT 0.090 1126.460 1241.940 1128.660 ;
        RECT 0.090 1125.300 1237.700 1126.460 ;
        RECT 1241.300 1125.300 1241.940 1126.460 ;
        RECT 0.090 1116.380 1241.940 1125.300 ;
        RECT 0.090 1115.220 0.700 1116.380 ;
        RECT 4.300 1115.220 1241.940 1116.380 ;
        RECT 0.090 1113.020 1241.940 1115.220 ;
        RECT 0.090 1111.860 1237.700 1113.020 ;
        RECT 1241.300 1111.860 1241.940 1113.020 ;
        RECT 0.090 1106.300 1241.940 1111.860 ;
        RECT 0.090 1105.140 0.700 1106.300 ;
        RECT 4.300 1105.140 1241.940 1106.300 ;
        RECT 0.090 1099.580 1241.940 1105.140 ;
        RECT 0.090 1098.420 1237.700 1099.580 ;
        RECT 1241.300 1098.420 1241.940 1099.580 ;
        RECT 0.090 1092.860 1241.940 1098.420 ;
        RECT 0.090 1091.700 0.700 1092.860 ;
        RECT 4.300 1091.700 1241.940 1092.860 ;
        RECT 0.090 1089.500 1241.940 1091.700 ;
        RECT 0.090 1088.340 1237.700 1089.500 ;
        RECT 1241.300 1088.340 1241.940 1089.500 ;
        RECT 0.090 1079.420 1241.940 1088.340 ;
        RECT 0.090 1078.260 0.700 1079.420 ;
        RECT 4.300 1078.260 1241.940 1079.420 ;
        RECT 0.090 1076.060 1241.940 1078.260 ;
        RECT 0.090 1074.900 1237.700 1076.060 ;
        RECT 1241.300 1074.900 1241.940 1076.060 ;
        RECT 0.090 1069.340 1241.940 1074.900 ;
        RECT 0.090 1068.180 0.700 1069.340 ;
        RECT 4.300 1068.180 1241.940 1069.340 ;
        RECT 0.090 1065.980 1241.940 1068.180 ;
        RECT 0.090 1064.820 1237.700 1065.980 ;
        RECT 1241.300 1064.820 1241.940 1065.980 ;
        RECT 0.090 1055.900 1241.940 1064.820 ;
        RECT 0.090 1054.740 0.700 1055.900 ;
        RECT 4.300 1054.740 1241.940 1055.900 ;
        RECT 0.090 1052.540 1241.940 1054.740 ;
        RECT 0.090 1051.380 1237.700 1052.540 ;
        RECT 1241.300 1051.380 1241.940 1052.540 ;
        RECT 0.090 1045.820 1241.940 1051.380 ;
        RECT 0.090 1044.660 0.700 1045.820 ;
        RECT 4.300 1044.660 1241.940 1045.820 ;
        RECT 0.090 1039.100 1241.940 1044.660 ;
        RECT 0.090 1037.940 1237.700 1039.100 ;
        RECT 1241.300 1037.940 1241.940 1039.100 ;
        RECT 0.090 1032.380 1241.940 1037.940 ;
        RECT 0.090 1031.220 0.700 1032.380 ;
        RECT 4.300 1031.220 1241.940 1032.380 ;
        RECT 0.090 1029.020 1241.940 1031.220 ;
        RECT 0.090 1027.860 1237.700 1029.020 ;
        RECT 1241.300 1027.860 1241.940 1029.020 ;
        RECT 0.090 1018.940 1241.940 1027.860 ;
        RECT 0.090 1017.780 0.700 1018.940 ;
        RECT 4.300 1017.780 1241.940 1018.940 ;
        RECT 0.090 1015.580 1241.940 1017.780 ;
        RECT 0.090 1014.420 1237.700 1015.580 ;
        RECT 1241.300 1014.420 1241.940 1015.580 ;
        RECT 0.090 1008.860 1241.940 1014.420 ;
        RECT 0.090 1007.700 0.700 1008.860 ;
        RECT 4.300 1007.700 1241.940 1008.860 ;
        RECT 0.090 1005.500 1241.940 1007.700 ;
        RECT 0.090 1004.340 1237.700 1005.500 ;
        RECT 1241.300 1004.340 1241.940 1005.500 ;
        RECT 0.090 995.420 1241.940 1004.340 ;
        RECT 0.090 994.260 0.700 995.420 ;
        RECT 4.300 994.260 1241.940 995.420 ;
        RECT 0.090 992.060 1241.940 994.260 ;
        RECT 0.090 990.900 1237.700 992.060 ;
        RECT 1241.300 990.900 1241.940 992.060 ;
        RECT 0.090 981.980 1241.940 990.900 ;
        RECT 0.090 980.820 0.700 981.980 ;
        RECT 4.300 980.820 1241.940 981.980 ;
        RECT 0.090 978.620 1241.940 980.820 ;
        RECT 0.090 977.460 1237.700 978.620 ;
        RECT 1241.300 977.460 1241.940 978.620 ;
        RECT 0.090 971.900 1241.940 977.460 ;
        RECT 0.090 970.740 0.700 971.900 ;
        RECT 4.300 970.740 1241.940 971.900 ;
        RECT 0.090 968.540 1241.940 970.740 ;
        RECT 0.090 967.380 1237.700 968.540 ;
        RECT 1241.300 967.380 1241.940 968.540 ;
        RECT 0.090 958.460 1241.940 967.380 ;
        RECT 0.090 957.300 0.700 958.460 ;
        RECT 4.300 957.300 1241.940 958.460 ;
        RECT 0.090 955.100 1241.940 957.300 ;
        RECT 0.090 953.940 1237.700 955.100 ;
        RECT 1241.300 953.940 1241.940 955.100 ;
        RECT 0.090 948.380 1241.940 953.940 ;
        RECT 0.090 947.220 0.700 948.380 ;
        RECT 4.300 947.220 1241.940 948.380 ;
        RECT 0.090 941.660 1241.940 947.220 ;
        RECT 0.090 940.500 1237.700 941.660 ;
        RECT 1241.300 940.500 1241.940 941.660 ;
        RECT 0.090 934.940 1241.940 940.500 ;
        RECT 0.090 933.780 0.700 934.940 ;
        RECT 4.300 933.780 1241.940 934.940 ;
        RECT 0.090 931.580 1241.940 933.780 ;
        RECT 0.090 930.420 1237.700 931.580 ;
        RECT 1241.300 930.420 1241.940 931.580 ;
        RECT 0.090 921.500 1241.940 930.420 ;
        RECT 0.090 920.340 0.700 921.500 ;
        RECT 4.300 920.340 1241.940 921.500 ;
        RECT 0.090 918.140 1241.940 920.340 ;
        RECT 0.090 916.980 1237.700 918.140 ;
        RECT 1241.300 916.980 1241.940 918.140 ;
        RECT 0.090 911.420 1241.940 916.980 ;
        RECT 0.090 910.260 0.700 911.420 ;
        RECT 4.300 910.260 1241.940 911.420 ;
        RECT 0.090 908.060 1241.940 910.260 ;
        RECT 0.090 906.900 1237.700 908.060 ;
        RECT 1241.300 906.900 1241.940 908.060 ;
        RECT 0.090 897.980 1241.940 906.900 ;
        RECT 0.090 896.820 0.700 897.980 ;
        RECT 4.300 896.820 1241.940 897.980 ;
        RECT 0.090 894.620 1241.940 896.820 ;
        RECT 0.090 893.460 1237.700 894.620 ;
        RECT 1241.300 893.460 1241.940 894.620 ;
        RECT 0.090 887.900 1241.940 893.460 ;
        RECT 0.090 886.740 0.700 887.900 ;
        RECT 4.300 886.740 1241.940 887.900 ;
        RECT 0.090 881.180 1241.940 886.740 ;
        RECT 0.090 880.020 1237.700 881.180 ;
        RECT 1241.300 880.020 1241.940 881.180 ;
        RECT 0.090 874.460 1241.940 880.020 ;
        RECT 0.090 873.300 0.700 874.460 ;
        RECT 4.300 873.300 1241.940 874.460 ;
        RECT 0.090 871.100 1241.940 873.300 ;
        RECT 0.090 869.940 1237.700 871.100 ;
        RECT 1241.300 869.940 1241.940 871.100 ;
        RECT 0.090 861.020 1241.940 869.940 ;
        RECT 0.090 859.860 0.700 861.020 ;
        RECT 4.300 859.860 1241.940 861.020 ;
        RECT 0.090 857.660 1241.940 859.860 ;
        RECT 0.090 856.500 1237.700 857.660 ;
        RECT 1241.300 856.500 1241.940 857.660 ;
        RECT 0.090 850.940 1241.940 856.500 ;
        RECT 0.090 849.780 0.700 850.940 ;
        RECT 4.300 849.780 1241.940 850.940 ;
        RECT 0.090 847.580 1241.940 849.780 ;
        RECT 0.090 846.420 1237.700 847.580 ;
        RECT 1241.300 846.420 1241.940 847.580 ;
        RECT 0.090 837.500 1241.940 846.420 ;
        RECT 0.090 836.340 0.700 837.500 ;
        RECT 4.300 836.340 1241.940 837.500 ;
        RECT 0.090 834.140 1241.940 836.340 ;
        RECT 0.090 832.980 1237.700 834.140 ;
        RECT 1241.300 832.980 1241.940 834.140 ;
        RECT 0.090 824.060 1241.940 832.980 ;
        RECT 0.090 822.900 0.700 824.060 ;
        RECT 4.300 822.900 1241.940 824.060 ;
        RECT 0.090 820.700 1241.940 822.900 ;
        RECT 0.090 819.540 1237.700 820.700 ;
        RECT 1241.300 819.540 1241.940 820.700 ;
        RECT 0.090 813.980 1241.940 819.540 ;
        RECT 0.090 812.820 0.700 813.980 ;
        RECT 4.300 812.820 1241.940 813.980 ;
        RECT 0.090 810.620 1241.940 812.820 ;
        RECT 0.090 809.460 1237.700 810.620 ;
        RECT 1241.300 809.460 1241.940 810.620 ;
        RECT 0.090 800.540 1241.940 809.460 ;
        RECT 0.090 799.380 0.700 800.540 ;
        RECT 4.300 799.380 1241.940 800.540 ;
        RECT 0.090 797.180 1241.940 799.380 ;
        RECT 0.090 796.020 1237.700 797.180 ;
        RECT 1241.300 796.020 1241.940 797.180 ;
        RECT 0.090 790.460 1241.940 796.020 ;
        RECT 0.090 789.300 0.700 790.460 ;
        RECT 4.300 789.300 1241.940 790.460 ;
        RECT 0.090 783.740 1241.940 789.300 ;
        RECT 0.090 782.580 1237.700 783.740 ;
        RECT 1241.300 782.580 1241.940 783.740 ;
        RECT 0.090 777.020 1241.940 782.580 ;
        RECT 0.090 775.860 0.700 777.020 ;
        RECT 4.300 775.860 1241.940 777.020 ;
        RECT 0.090 773.660 1241.940 775.860 ;
        RECT 0.090 772.500 1237.700 773.660 ;
        RECT 1241.300 772.500 1241.940 773.660 ;
        RECT 0.090 763.580 1241.940 772.500 ;
        RECT 0.090 762.420 0.700 763.580 ;
        RECT 4.300 762.420 1241.940 763.580 ;
        RECT 0.090 760.220 1241.940 762.420 ;
        RECT 0.090 759.060 1237.700 760.220 ;
        RECT 1241.300 759.060 1241.940 760.220 ;
        RECT 0.090 753.500 1241.940 759.060 ;
        RECT 0.090 752.340 0.700 753.500 ;
        RECT 4.300 752.340 1241.940 753.500 ;
        RECT 0.090 750.140 1241.940 752.340 ;
        RECT 0.090 748.980 1237.700 750.140 ;
        RECT 1241.300 748.980 1241.940 750.140 ;
        RECT 0.090 740.060 1241.940 748.980 ;
        RECT 0.090 738.900 0.700 740.060 ;
        RECT 4.300 738.900 1241.940 740.060 ;
        RECT 0.090 736.700 1241.940 738.900 ;
        RECT 0.090 735.540 1237.700 736.700 ;
        RECT 1241.300 735.540 1241.940 736.700 ;
        RECT 0.090 726.620 1241.940 735.540 ;
        RECT 0.090 725.460 0.700 726.620 ;
        RECT 4.300 725.460 1241.940 726.620 ;
        RECT 0.090 723.260 1241.940 725.460 ;
        RECT 0.090 722.100 1237.700 723.260 ;
        RECT 1241.300 722.100 1241.940 723.260 ;
        RECT 0.090 716.540 1241.940 722.100 ;
        RECT 0.090 715.380 0.700 716.540 ;
        RECT 4.300 715.380 1241.940 716.540 ;
        RECT 0.090 713.180 1241.940 715.380 ;
        RECT 0.090 712.020 1237.700 713.180 ;
        RECT 1241.300 712.020 1241.940 713.180 ;
        RECT 0.090 703.100 1241.940 712.020 ;
        RECT 0.090 701.940 0.700 703.100 ;
        RECT 4.300 701.940 1241.940 703.100 ;
        RECT 0.090 699.740 1241.940 701.940 ;
        RECT 0.090 698.580 1237.700 699.740 ;
        RECT 1241.300 698.580 1241.940 699.740 ;
        RECT 0.090 693.020 1241.940 698.580 ;
        RECT 0.090 691.860 0.700 693.020 ;
        RECT 4.300 691.860 1241.940 693.020 ;
        RECT 0.090 689.660 1241.940 691.860 ;
        RECT 0.090 688.500 1237.700 689.660 ;
        RECT 1241.300 688.500 1241.940 689.660 ;
        RECT 0.090 679.580 1241.940 688.500 ;
        RECT 0.090 678.420 0.700 679.580 ;
        RECT 4.300 678.420 1241.940 679.580 ;
        RECT 0.090 676.220 1241.940 678.420 ;
        RECT 0.090 675.060 1237.700 676.220 ;
        RECT 1241.300 675.060 1241.940 676.220 ;
        RECT 0.090 666.140 1241.940 675.060 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 1241.940 666.140 ;
        RECT 0.090 662.780 1241.940 664.980 ;
        RECT 0.090 661.620 1237.700 662.780 ;
        RECT 1241.300 661.620 1241.940 662.780 ;
        RECT 0.090 656.060 1241.940 661.620 ;
        RECT 0.090 654.900 0.700 656.060 ;
        RECT 4.300 654.900 1241.940 656.060 ;
        RECT 0.090 652.700 1241.940 654.900 ;
        RECT 0.090 651.540 1237.700 652.700 ;
        RECT 1241.300 651.540 1241.940 652.700 ;
        RECT 0.090 642.620 1241.940 651.540 ;
        RECT 0.090 641.460 0.700 642.620 ;
        RECT 4.300 641.460 1241.940 642.620 ;
        RECT 0.090 639.260 1241.940 641.460 ;
        RECT 0.090 638.100 1237.700 639.260 ;
        RECT 1241.300 638.100 1241.940 639.260 ;
        RECT 0.090 632.540 1241.940 638.100 ;
        RECT 0.090 631.380 0.700 632.540 ;
        RECT 4.300 631.380 1241.940 632.540 ;
        RECT 0.090 625.820 1241.940 631.380 ;
        RECT 0.090 624.660 1237.700 625.820 ;
        RECT 1241.300 624.660 1241.940 625.820 ;
        RECT 0.090 619.100 1241.940 624.660 ;
        RECT 0.090 617.940 0.700 619.100 ;
        RECT 4.300 617.940 1241.940 619.100 ;
        RECT 0.090 615.740 1241.940 617.940 ;
        RECT 0.090 614.580 1237.700 615.740 ;
        RECT 1241.300 614.580 1241.940 615.740 ;
        RECT 0.090 605.660 1241.940 614.580 ;
        RECT 0.090 604.500 0.700 605.660 ;
        RECT 4.300 604.500 1241.940 605.660 ;
        RECT 0.090 602.300 1241.940 604.500 ;
        RECT 0.090 601.140 1237.700 602.300 ;
        RECT 1241.300 601.140 1241.940 602.300 ;
        RECT 0.090 595.580 1241.940 601.140 ;
        RECT 0.090 594.420 0.700 595.580 ;
        RECT 4.300 594.420 1241.940 595.580 ;
        RECT 0.090 592.220 1241.940 594.420 ;
        RECT 0.090 591.060 1237.700 592.220 ;
        RECT 1241.300 591.060 1241.940 592.220 ;
        RECT 0.090 582.140 1241.940 591.060 ;
        RECT 0.090 580.980 0.700 582.140 ;
        RECT 4.300 580.980 1241.940 582.140 ;
        RECT 0.090 578.780 1241.940 580.980 ;
        RECT 0.090 577.620 1237.700 578.780 ;
        RECT 1241.300 577.620 1241.940 578.780 ;
        RECT 0.090 568.700 1241.940 577.620 ;
        RECT 0.090 567.540 0.700 568.700 ;
        RECT 4.300 567.540 1241.940 568.700 ;
        RECT 0.090 565.340 1241.940 567.540 ;
        RECT 0.090 564.180 1237.700 565.340 ;
        RECT 1241.300 564.180 1241.940 565.340 ;
        RECT 0.090 558.620 1241.940 564.180 ;
        RECT 0.090 557.460 0.700 558.620 ;
        RECT 4.300 557.460 1241.940 558.620 ;
        RECT 0.090 555.260 1241.940 557.460 ;
        RECT 0.090 554.100 1237.700 555.260 ;
        RECT 1241.300 554.100 1241.940 555.260 ;
        RECT 0.090 545.180 1241.940 554.100 ;
        RECT 0.090 544.020 0.700 545.180 ;
        RECT 4.300 544.020 1241.940 545.180 ;
        RECT 0.090 541.820 1241.940 544.020 ;
        RECT 0.090 540.660 1237.700 541.820 ;
        RECT 1241.300 540.660 1241.940 541.820 ;
        RECT 0.090 535.100 1241.940 540.660 ;
        RECT 0.090 533.940 0.700 535.100 ;
        RECT 4.300 533.940 1241.940 535.100 ;
        RECT 0.090 531.740 1241.940 533.940 ;
        RECT 0.090 530.580 1237.700 531.740 ;
        RECT 1241.300 530.580 1241.940 531.740 ;
        RECT 0.090 521.660 1241.940 530.580 ;
        RECT 0.090 520.500 0.700 521.660 ;
        RECT 4.300 520.500 1241.940 521.660 ;
        RECT 0.090 518.300 1241.940 520.500 ;
        RECT 0.090 517.140 1237.700 518.300 ;
        RECT 1241.300 517.140 1241.940 518.300 ;
        RECT 0.090 508.220 1241.940 517.140 ;
        RECT 0.090 507.060 0.700 508.220 ;
        RECT 4.300 507.060 1241.940 508.220 ;
        RECT 0.090 504.860 1241.940 507.060 ;
        RECT 0.090 503.700 1237.700 504.860 ;
        RECT 1241.300 503.700 1241.940 504.860 ;
        RECT 0.090 498.140 1241.940 503.700 ;
        RECT 0.090 496.980 0.700 498.140 ;
        RECT 4.300 496.980 1241.940 498.140 ;
        RECT 0.090 494.780 1241.940 496.980 ;
        RECT 0.090 493.620 1237.700 494.780 ;
        RECT 1241.300 493.620 1241.940 494.780 ;
        RECT 0.090 484.700 1241.940 493.620 ;
        RECT 0.090 483.540 0.700 484.700 ;
        RECT 4.300 483.540 1241.940 484.700 ;
        RECT 0.090 481.340 1241.940 483.540 ;
        RECT 0.090 480.180 1237.700 481.340 ;
        RECT 1241.300 480.180 1241.940 481.340 ;
        RECT 0.090 474.620 1241.940 480.180 ;
        RECT 0.090 473.460 0.700 474.620 ;
        RECT 4.300 473.460 1241.940 474.620 ;
        RECT 0.090 467.900 1241.940 473.460 ;
        RECT 0.090 466.740 1237.700 467.900 ;
        RECT 1241.300 466.740 1241.940 467.900 ;
        RECT 0.090 461.180 1241.940 466.740 ;
        RECT 0.090 460.020 0.700 461.180 ;
        RECT 4.300 460.020 1241.940 461.180 ;
        RECT 0.090 457.820 1241.940 460.020 ;
        RECT 0.090 456.660 1237.700 457.820 ;
        RECT 1241.300 456.660 1241.940 457.820 ;
        RECT 0.090 447.740 1241.940 456.660 ;
        RECT 0.090 446.580 0.700 447.740 ;
        RECT 4.300 446.580 1241.940 447.740 ;
        RECT 0.090 444.380 1241.940 446.580 ;
        RECT 0.090 443.220 1237.700 444.380 ;
        RECT 1241.300 443.220 1241.940 444.380 ;
        RECT 0.090 437.660 1241.940 443.220 ;
        RECT 0.090 436.500 0.700 437.660 ;
        RECT 4.300 436.500 1241.940 437.660 ;
        RECT 0.090 434.300 1241.940 436.500 ;
        RECT 0.090 433.140 1237.700 434.300 ;
        RECT 1241.300 433.140 1241.940 434.300 ;
        RECT 0.090 424.220 1241.940 433.140 ;
        RECT 0.090 423.060 0.700 424.220 ;
        RECT 4.300 423.060 1241.940 424.220 ;
        RECT 0.090 420.860 1241.940 423.060 ;
        RECT 0.090 419.700 1237.700 420.860 ;
        RECT 1241.300 419.700 1241.940 420.860 ;
        RECT 0.090 410.780 1241.940 419.700 ;
        RECT 0.090 409.620 0.700 410.780 ;
        RECT 4.300 409.620 1241.940 410.780 ;
        RECT 0.090 407.420 1241.940 409.620 ;
        RECT 0.090 406.260 1237.700 407.420 ;
        RECT 1241.300 406.260 1241.940 407.420 ;
        RECT 0.090 400.700 1241.940 406.260 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 1241.940 400.700 ;
        RECT 0.090 397.340 1241.940 399.540 ;
        RECT 0.090 396.180 1237.700 397.340 ;
        RECT 1241.300 396.180 1241.940 397.340 ;
        RECT 0.090 387.260 1241.940 396.180 ;
        RECT 0.090 386.100 0.700 387.260 ;
        RECT 4.300 386.100 1241.940 387.260 ;
        RECT 0.090 383.900 1241.940 386.100 ;
        RECT 0.090 382.740 1237.700 383.900 ;
        RECT 1241.300 382.740 1241.940 383.900 ;
        RECT 0.090 377.180 1241.940 382.740 ;
        RECT 0.090 376.020 0.700 377.180 ;
        RECT 4.300 376.020 1241.940 377.180 ;
        RECT 0.090 370.460 1241.940 376.020 ;
        RECT 0.090 369.300 1237.700 370.460 ;
        RECT 1241.300 369.300 1241.940 370.460 ;
        RECT 0.090 363.740 1241.940 369.300 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 1241.940 363.740 ;
        RECT 0.090 360.380 1241.940 362.580 ;
        RECT 0.090 359.220 1237.700 360.380 ;
        RECT 1241.300 359.220 1241.940 360.380 ;
        RECT 0.090 350.300 1241.940 359.220 ;
        RECT 0.090 349.140 0.700 350.300 ;
        RECT 4.300 349.140 1241.940 350.300 ;
        RECT 0.090 346.940 1241.940 349.140 ;
        RECT 0.090 345.780 1237.700 346.940 ;
        RECT 1241.300 345.780 1241.940 346.940 ;
        RECT 0.090 340.220 1241.940 345.780 ;
        RECT 0.090 339.060 0.700 340.220 ;
        RECT 4.300 339.060 1241.940 340.220 ;
        RECT 0.090 336.860 1241.940 339.060 ;
        RECT 0.090 335.700 1237.700 336.860 ;
        RECT 1241.300 335.700 1241.940 336.860 ;
        RECT 0.090 326.780 1241.940 335.700 ;
        RECT 0.090 325.620 0.700 326.780 ;
        RECT 4.300 325.620 1241.940 326.780 ;
        RECT 0.090 323.420 1241.940 325.620 ;
        RECT 0.090 322.260 1237.700 323.420 ;
        RECT 1241.300 322.260 1241.940 323.420 ;
        RECT 0.090 316.700 1241.940 322.260 ;
        RECT 0.090 315.540 0.700 316.700 ;
        RECT 4.300 315.540 1241.940 316.700 ;
        RECT 0.090 309.980 1241.940 315.540 ;
        RECT 0.090 308.820 1237.700 309.980 ;
        RECT 1241.300 308.820 1241.940 309.980 ;
        RECT 0.090 303.260 1241.940 308.820 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 1241.940 303.260 ;
        RECT 0.090 299.900 1241.940 302.100 ;
        RECT 0.090 298.740 1237.700 299.900 ;
        RECT 1241.300 298.740 1241.940 299.900 ;
        RECT 0.090 289.820 1241.940 298.740 ;
        RECT 0.090 288.660 0.700 289.820 ;
        RECT 4.300 288.660 1241.940 289.820 ;
        RECT 0.090 286.460 1241.940 288.660 ;
        RECT 0.090 285.300 1237.700 286.460 ;
        RECT 1241.300 285.300 1241.940 286.460 ;
        RECT 0.090 279.740 1241.940 285.300 ;
        RECT 0.090 278.580 0.700 279.740 ;
        RECT 4.300 278.580 1241.940 279.740 ;
        RECT 0.090 276.380 1241.940 278.580 ;
        RECT 0.090 275.220 1237.700 276.380 ;
        RECT 1241.300 275.220 1241.940 276.380 ;
        RECT 0.090 266.300 1241.940 275.220 ;
        RECT 0.090 265.140 0.700 266.300 ;
        RECT 4.300 265.140 1241.940 266.300 ;
        RECT 0.090 262.940 1241.940 265.140 ;
        RECT 0.090 261.780 1237.700 262.940 ;
        RECT 1241.300 261.780 1241.940 262.940 ;
        RECT 0.090 252.860 1241.940 261.780 ;
        RECT 0.090 251.700 0.700 252.860 ;
        RECT 4.300 251.700 1241.940 252.860 ;
        RECT 0.090 249.500 1241.940 251.700 ;
        RECT 0.090 248.340 1237.700 249.500 ;
        RECT 1241.300 248.340 1241.940 249.500 ;
        RECT 0.090 242.780 1241.940 248.340 ;
        RECT 0.090 241.620 0.700 242.780 ;
        RECT 4.300 241.620 1241.940 242.780 ;
        RECT 0.090 239.420 1241.940 241.620 ;
        RECT 0.090 238.260 1237.700 239.420 ;
        RECT 1241.300 238.260 1241.940 239.420 ;
        RECT 0.090 229.340 1241.940 238.260 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 1241.940 229.340 ;
        RECT 0.090 225.980 1241.940 228.180 ;
        RECT 0.090 224.820 1237.700 225.980 ;
        RECT 1241.300 224.820 1241.940 225.980 ;
        RECT 0.090 219.260 1241.940 224.820 ;
        RECT 0.090 218.100 0.700 219.260 ;
        RECT 4.300 218.100 1241.940 219.260 ;
        RECT 0.090 212.540 1241.940 218.100 ;
        RECT 0.090 211.380 1237.700 212.540 ;
        RECT 1241.300 211.380 1241.940 212.540 ;
        RECT 0.090 205.820 1241.940 211.380 ;
        RECT 0.090 204.660 0.700 205.820 ;
        RECT 4.300 204.660 1241.940 205.820 ;
        RECT 0.090 202.460 1241.940 204.660 ;
        RECT 0.090 201.300 1237.700 202.460 ;
        RECT 1241.300 201.300 1241.940 202.460 ;
        RECT 0.090 192.380 1241.940 201.300 ;
        RECT 0.090 191.220 0.700 192.380 ;
        RECT 4.300 191.220 1241.940 192.380 ;
        RECT 0.090 189.020 1241.940 191.220 ;
        RECT 0.090 187.860 1237.700 189.020 ;
        RECT 1241.300 187.860 1241.940 189.020 ;
        RECT 0.090 182.300 1241.940 187.860 ;
        RECT 0.090 181.140 0.700 182.300 ;
        RECT 4.300 181.140 1241.940 182.300 ;
        RECT 0.090 178.940 1241.940 181.140 ;
        RECT 0.090 177.780 1237.700 178.940 ;
        RECT 1241.300 177.780 1241.940 178.940 ;
        RECT 0.090 168.860 1241.940 177.780 ;
        RECT 0.090 167.700 0.700 168.860 ;
        RECT 4.300 167.700 1241.940 168.860 ;
        RECT 0.090 165.500 1241.940 167.700 ;
        RECT 0.090 164.340 1237.700 165.500 ;
        RECT 1241.300 164.340 1241.940 165.500 ;
        RECT 0.090 158.780 1241.940 164.340 ;
        RECT 0.090 157.620 0.700 158.780 ;
        RECT 4.300 157.620 1241.940 158.780 ;
        RECT 0.090 152.060 1241.940 157.620 ;
        RECT 0.090 150.900 1237.700 152.060 ;
        RECT 1241.300 150.900 1241.940 152.060 ;
        RECT 0.090 145.340 1241.940 150.900 ;
        RECT 0.090 144.180 0.700 145.340 ;
        RECT 4.300 144.180 1241.940 145.340 ;
        RECT 0.090 141.980 1241.940 144.180 ;
        RECT 0.090 140.820 1237.700 141.980 ;
        RECT 1241.300 140.820 1241.940 141.980 ;
        RECT 0.090 131.900 1241.940 140.820 ;
        RECT 0.090 130.740 0.700 131.900 ;
        RECT 4.300 130.740 1241.940 131.900 ;
        RECT 0.090 128.540 1241.940 130.740 ;
        RECT 0.090 127.380 1237.700 128.540 ;
        RECT 1241.300 127.380 1241.940 128.540 ;
        RECT 0.090 121.820 1241.940 127.380 ;
        RECT 0.090 120.660 0.700 121.820 ;
        RECT 4.300 120.660 1241.940 121.820 ;
        RECT 0.090 118.460 1241.940 120.660 ;
        RECT 0.090 117.300 1237.700 118.460 ;
        RECT 1241.300 117.300 1241.940 118.460 ;
        RECT 0.090 108.380 1241.940 117.300 ;
        RECT 0.090 107.220 0.700 108.380 ;
        RECT 4.300 107.220 1241.940 108.380 ;
        RECT 0.090 105.020 1241.940 107.220 ;
        RECT 0.090 103.860 1237.700 105.020 ;
        RECT 1241.300 103.860 1241.940 105.020 ;
        RECT 0.090 94.940 1241.940 103.860 ;
        RECT 0.090 93.780 0.700 94.940 ;
        RECT 4.300 93.780 1241.940 94.940 ;
        RECT 0.090 91.580 1241.940 93.780 ;
        RECT 0.090 90.420 1237.700 91.580 ;
        RECT 1241.300 90.420 1241.940 91.580 ;
        RECT 0.090 84.860 1241.940 90.420 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 1241.940 84.860 ;
        RECT 0.090 81.500 1241.940 83.700 ;
        RECT 0.090 80.340 1237.700 81.500 ;
        RECT 1241.300 80.340 1241.940 81.500 ;
        RECT 0.090 71.420 1241.940 80.340 ;
        RECT 0.090 70.260 0.700 71.420 ;
        RECT 4.300 70.260 1241.940 71.420 ;
        RECT 0.090 68.060 1241.940 70.260 ;
        RECT 0.090 66.900 1237.700 68.060 ;
        RECT 1241.300 66.900 1241.940 68.060 ;
        RECT 0.090 61.340 1241.940 66.900 ;
        RECT 0.090 60.180 0.700 61.340 ;
        RECT 4.300 60.180 1241.940 61.340 ;
        RECT 0.090 54.620 1241.940 60.180 ;
        RECT 0.090 53.460 1237.700 54.620 ;
        RECT 1241.300 53.460 1241.940 54.620 ;
        RECT 0.090 47.900 1241.940 53.460 ;
        RECT 0.090 46.740 0.700 47.900 ;
        RECT 4.300 46.740 1241.940 47.900 ;
        RECT 0.090 44.540 1241.940 46.740 ;
        RECT 0.090 43.380 1237.700 44.540 ;
        RECT 1241.300 43.380 1241.940 44.540 ;
        RECT 0.090 34.460 1241.940 43.380 ;
        RECT 0.090 33.300 0.700 34.460 ;
        RECT 4.300 33.300 1241.940 34.460 ;
        RECT 0.090 31.100 1241.940 33.300 ;
        RECT 0.090 29.940 1237.700 31.100 ;
        RECT 1241.300 29.940 1241.940 31.100 ;
        RECT 0.090 24.380 1241.940 29.940 ;
        RECT 0.090 23.220 0.700 24.380 ;
        RECT 4.300 23.220 1241.940 24.380 ;
        RECT 0.090 21.020 1241.940 23.220 ;
        RECT 0.090 19.860 1237.700 21.020 ;
        RECT 1241.300 19.860 1241.940 21.020 ;
        RECT 0.090 10.940 1241.940 19.860 ;
        RECT 0.090 9.780 0.700 10.940 ;
        RECT 4.300 9.780 1241.940 10.940 ;
        RECT 0.090 7.980 1241.940 9.780 ;
      LAYER Metal4 ;
        RECT 21.420 15.080 21.940 1240.870 ;
        RECT 24.140 15.080 98.740 1240.870 ;
        RECT 100.940 15.080 175.540 1240.870 ;
        RECT 177.740 15.080 252.340 1240.870 ;
        RECT 254.540 15.080 329.140 1240.870 ;
        RECT 331.340 15.080 405.940 1240.870 ;
        RECT 408.140 15.080 482.740 1240.870 ;
        RECT 484.940 15.080 559.540 1240.870 ;
        RECT 561.740 15.080 636.340 1240.870 ;
        RECT 638.540 15.080 713.140 1240.870 ;
        RECT 715.340 15.080 789.940 1240.870 ;
        RECT 792.140 15.080 866.740 1240.870 ;
        RECT 868.940 15.080 943.540 1240.870 ;
        RECT 945.740 15.080 1020.340 1240.870 ;
        RECT 1022.540 15.080 1097.140 1240.870 ;
        RECT 1099.340 15.080 1173.940 1240.870 ;
        RECT 1176.140 15.080 1226.260 1240.870 ;
        RECT 21.420 13.530 1226.260 15.080 ;
  END
END aes_core
END LIBRARY

