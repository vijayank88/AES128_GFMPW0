magic
tech gf180mcuC
magscale 1 5
timestamp 1670062326
<< obsm1 >>
rect 672 855 123480 124294
<< metal2 >>
rect 336 125592 392 125892
rect 1344 125592 1400 125892
rect 2688 125592 2744 125892
rect 3696 125592 3752 125892
rect 5040 125592 5096 125892
rect 6384 125592 6440 125892
rect 7392 125592 7448 125892
rect 8736 125592 8792 125892
rect 10080 125592 10136 125892
rect 11088 125592 11144 125892
rect 12432 125592 12488 125892
rect 13440 125592 13496 125892
rect 14784 125592 14840 125892
rect 16128 125592 16184 125892
rect 17136 125592 17192 125892
rect 18480 125592 18536 125892
rect 19488 125592 19544 125892
rect 20832 125592 20888 125892
rect 22176 125592 22232 125892
rect 23184 125592 23240 125892
rect 24528 125592 24584 125892
rect 25872 125592 25928 125892
rect 26880 125592 26936 125892
rect 28224 125592 28280 125892
rect 29232 125592 29288 125892
rect 30576 125592 30632 125892
rect 31920 125592 31976 125892
rect 32928 125592 32984 125892
rect 34272 125592 34328 125892
rect 35280 125592 35336 125892
rect 36624 125592 36680 125892
rect 37968 125592 38024 125892
rect 38976 125592 39032 125892
rect 40320 125592 40376 125892
rect 41664 125592 41720 125892
rect 42672 125592 42728 125892
rect 44016 125592 44072 125892
rect 45024 125592 45080 125892
rect 46368 125592 46424 125892
rect 47712 125592 47768 125892
rect 48720 125592 48776 125892
rect 50064 125592 50120 125892
rect 51408 125592 51464 125892
rect 52416 125592 52472 125892
rect 53760 125592 53816 125892
rect 54768 125592 54824 125892
rect 56112 125592 56168 125892
rect 57456 125592 57512 125892
rect 58464 125592 58520 125892
rect 59808 125592 59864 125892
rect 60816 125592 60872 125892
rect 62160 125592 62216 125892
rect 63504 125592 63560 125892
rect 64512 125592 64568 125892
rect 65856 125592 65912 125892
rect 67200 125592 67256 125892
rect 68208 125592 68264 125892
rect 69552 125592 69608 125892
rect 70560 125592 70616 125892
rect 71904 125592 71960 125892
rect 73248 125592 73304 125892
rect 74256 125592 74312 125892
rect 75600 125592 75656 125892
rect 76608 125592 76664 125892
rect 77952 125592 78008 125892
rect 79296 125592 79352 125892
rect 80304 125592 80360 125892
rect 81648 125592 81704 125892
rect 82992 125592 83048 125892
rect 84000 125592 84056 125892
rect 85344 125592 85400 125892
rect 86352 125592 86408 125892
rect 87696 125592 87752 125892
rect 89040 125592 89096 125892
rect 90048 125592 90104 125892
rect 91392 125592 91448 125892
rect 92400 125592 92456 125892
rect 93744 125592 93800 125892
rect 95088 125592 95144 125892
rect 96096 125592 96152 125892
rect 97440 125592 97496 125892
rect 98784 125592 98840 125892
rect 99792 125592 99848 125892
rect 101136 125592 101192 125892
rect 102144 125592 102200 125892
rect 103488 125592 103544 125892
rect 104832 125592 104888 125892
rect 105840 125592 105896 125892
rect 107184 125592 107240 125892
rect 108192 125592 108248 125892
rect 109536 125592 109592 125892
rect 110880 125592 110936 125892
rect 111888 125592 111944 125892
rect 113232 125592 113288 125892
rect 114576 125592 114632 125892
rect 115584 125592 115640 125892
rect 116928 125592 116984 125892
rect 117936 125592 117992 125892
rect 119280 125592 119336 125892
rect 120624 125592 120680 125892
rect 121632 125592 121688 125892
rect 122976 125592 123032 125892
rect 123984 125592 124040 125892
rect 0 100 56 400
rect 1008 100 1064 400
rect 2352 100 2408 400
rect 3360 100 3416 400
rect 4704 100 4760 400
rect 6048 100 6104 400
rect 7056 100 7112 400
rect 8400 100 8456 400
rect 9408 100 9464 400
rect 10752 100 10808 400
rect 12096 100 12152 400
rect 13104 100 13160 400
rect 14448 100 14504 400
rect 15792 100 15848 400
rect 16800 100 16856 400
rect 18144 100 18200 400
rect 19152 100 19208 400
rect 20496 100 20552 400
rect 21840 100 21896 400
rect 22848 100 22904 400
rect 24192 100 24248 400
rect 25200 100 25256 400
rect 26544 100 26600 400
rect 27888 100 27944 400
rect 28896 100 28952 400
rect 30240 100 30296 400
rect 31584 100 31640 400
rect 32592 100 32648 400
rect 33936 100 33992 400
rect 34944 100 35000 400
rect 36288 100 36344 400
rect 37632 100 37688 400
rect 38640 100 38696 400
rect 39984 100 40040 400
rect 40992 100 41048 400
rect 42336 100 42392 400
rect 43680 100 43736 400
rect 44688 100 44744 400
rect 46032 100 46088 400
rect 47376 100 47432 400
rect 48384 100 48440 400
rect 49728 100 49784 400
rect 50736 100 50792 400
rect 52080 100 52136 400
rect 53424 100 53480 400
rect 54432 100 54488 400
rect 55776 100 55832 400
rect 56784 100 56840 400
rect 58128 100 58184 400
rect 59472 100 59528 400
rect 60480 100 60536 400
rect 61824 100 61880 400
rect 63168 100 63224 400
rect 64176 100 64232 400
rect 65520 100 65576 400
rect 66528 100 66584 400
rect 67872 100 67928 400
rect 69216 100 69272 400
rect 70224 100 70280 400
rect 71568 100 71624 400
rect 72576 100 72632 400
rect 73920 100 73976 400
rect 75264 100 75320 400
rect 76272 100 76328 400
rect 77616 100 77672 400
rect 78960 100 79016 400
rect 79968 100 80024 400
rect 81312 100 81368 400
rect 82320 100 82376 400
rect 83664 100 83720 400
rect 85008 100 85064 400
rect 86016 100 86072 400
rect 87360 100 87416 400
rect 88704 100 88760 400
rect 89712 100 89768 400
rect 91056 100 91112 400
rect 92064 100 92120 400
rect 93408 100 93464 400
rect 94752 100 94808 400
rect 95760 100 95816 400
rect 97104 100 97160 400
rect 98112 100 98168 400
rect 99456 100 99512 400
rect 100800 100 100856 400
rect 101808 100 101864 400
rect 103152 100 103208 400
rect 104496 100 104552 400
rect 105504 100 105560 400
rect 106848 100 106904 400
rect 107856 100 107912 400
rect 109200 100 109256 400
rect 110544 100 110600 400
rect 111552 100 111608 400
rect 112896 100 112952 400
rect 113904 100 113960 400
rect 115248 100 115304 400
rect 116592 100 116648 400
rect 117600 100 117656 400
rect 118944 100 119000 400
rect 120288 100 120344 400
rect 121296 100 121352 400
rect 122640 100 122696 400
rect 123648 100 123704 400
<< obsm2 >>
rect 14 125562 306 125650
rect 422 125562 1314 125650
rect 1430 125562 2658 125650
rect 2774 125562 3666 125650
rect 3782 125562 5010 125650
rect 5126 125562 6354 125650
rect 6470 125562 7362 125650
rect 7478 125562 8706 125650
rect 8822 125562 10050 125650
rect 10166 125562 11058 125650
rect 11174 125562 12402 125650
rect 12518 125562 13410 125650
rect 13526 125562 14754 125650
rect 14870 125562 16098 125650
rect 16214 125562 17106 125650
rect 17222 125562 18450 125650
rect 18566 125562 19458 125650
rect 19574 125562 20802 125650
rect 20918 125562 22146 125650
rect 22262 125562 23154 125650
rect 23270 125562 24498 125650
rect 24614 125562 25842 125650
rect 25958 125562 26850 125650
rect 26966 125562 28194 125650
rect 28310 125562 29202 125650
rect 29318 125562 30546 125650
rect 30662 125562 31890 125650
rect 32006 125562 32898 125650
rect 33014 125562 34242 125650
rect 34358 125562 35250 125650
rect 35366 125562 36594 125650
rect 36710 125562 37938 125650
rect 38054 125562 38946 125650
rect 39062 125562 40290 125650
rect 40406 125562 41634 125650
rect 41750 125562 42642 125650
rect 42758 125562 43986 125650
rect 44102 125562 44994 125650
rect 45110 125562 46338 125650
rect 46454 125562 47682 125650
rect 47798 125562 48690 125650
rect 48806 125562 50034 125650
rect 50150 125562 51378 125650
rect 51494 125562 52386 125650
rect 52502 125562 53730 125650
rect 53846 125562 54738 125650
rect 54854 125562 56082 125650
rect 56198 125562 57426 125650
rect 57542 125562 58434 125650
rect 58550 125562 59778 125650
rect 59894 125562 60786 125650
rect 60902 125562 62130 125650
rect 62246 125562 63474 125650
rect 63590 125562 64482 125650
rect 64598 125562 65826 125650
rect 65942 125562 67170 125650
rect 67286 125562 68178 125650
rect 68294 125562 69522 125650
rect 69638 125562 70530 125650
rect 70646 125562 71874 125650
rect 71990 125562 73218 125650
rect 73334 125562 74226 125650
rect 74342 125562 75570 125650
rect 75686 125562 76578 125650
rect 76694 125562 77922 125650
rect 78038 125562 79266 125650
rect 79382 125562 80274 125650
rect 80390 125562 81618 125650
rect 81734 125562 82962 125650
rect 83078 125562 83970 125650
rect 84086 125562 85314 125650
rect 85430 125562 86322 125650
rect 86438 125562 87666 125650
rect 87782 125562 89010 125650
rect 89126 125562 90018 125650
rect 90134 125562 91362 125650
rect 91478 125562 92370 125650
rect 92486 125562 93714 125650
rect 93830 125562 95058 125650
rect 95174 125562 96066 125650
rect 96182 125562 97410 125650
rect 97526 125562 98754 125650
rect 98870 125562 99762 125650
rect 99878 125562 101106 125650
rect 101222 125562 102114 125650
rect 102230 125562 103458 125650
rect 103574 125562 104802 125650
rect 104918 125562 105810 125650
rect 105926 125562 107154 125650
rect 107270 125562 108162 125650
rect 108278 125562 109506 125650
rect 109622 125562 110850 125650
rect 110966 125562 111858 125650
rect 111974 125562 113202 125650
rect 113318 125562 114546 125650
rect 114662 125562 115554 125650
rect 115670 125562 116898 125650
rect 117014 125562 117906 125650
rect 118022 125562 119250 125650
rect 119366 125562 120594 125650
rect 120710 125562 121602 125650
rect 121718 125562 122946 125650
rect 123062 125562 123578 125650
rect 14 430 123578 125562
rect 86 400 978 430
rect 1094 400 2322 430
rect 2438 400 3330 430
rect 3446 400 4674 430
rect 4790 400 6018 430
rect 6134 400 7026 430
rect 7142 400 8370 430
rect 8486 400 9378 430
rect 9494 400 10722 430
rect 10838 400 12066 430
rect 12182 400 13074 430
rect 13190 400 14418 430
rect 14534 400 15762 430
rect 15878 400 16770 430
rect 16886 400 18114 430
rect 18230 400 19122 430
rect 19238 400 20466 430
rect 20582 400 21810 430
rect 21926 400 22818 430
rect 22934 400 24162 430
rect 24278 400 25170 430
rect 25286 400 26514 430
rect 26630 400 27858 430
rect 27974 400 28866 430
rect 28982 400 30210 430
rect 30326 400 31554 430
rect 31670 400 32562 430
rect 32678 400 33906 430
rect 34022 400 34914 430
rect 35030 400 36258 430
rect 36374 400 37602 430
rect 37718 400 38610 430
rect 38726 400 39954 430
rect 40070 400 40962 430
rect 41078 400 42306 430
rect 42422 400 43650 430
rect 43766 400 44658 430
rect 44774 400 46002 430
rect 46118 400 47346 430
rect 47462 400 48354 430
rect 48470 400 49698 430
rect 49814 400 50706 430
rect 50822 400 52050 430
rect 52166 400 53394 430
rect 53510 400 54402 430
rect 54518 400 55746 430
rect 55862 400 56754 430
rect 56870 400 58098 430
rect 58214 400 59442 430
rect 59558 400 60450 430
rect 60566 400 61794 430
rect 61910 400 63138 430
rect 63254 400 64146 430
rect 64262 400 65490 430
rect 65606 400 66498 430
rect 66614 400 67842 430
rect 67958 400 69186 430
rect 69302 400 70194 430
rect 70310 400 71538 430
rect 71654 400 72546 430
rect 72662 400 73890 430
rect 74006 400 75234 430
rect 75350 400 76242 430
rect 76358 400 77586 430
rect 77702 400 78930 430
rect 79046 400 79938 430
rect 80054 400 81282 430
rect 81398 400 82290 430
rect 82406 400 83634 430
rect 83750 400 84978 430
rect 85094 400 85986 430
rect 86102 400 87330 430
rect 87446 400 88674 430
rect 88790 400 89682 430
rect 89798 400 91026 430
rect 91142 400 92034 430
rect 92150 400 93378 430
rect 93494 400 94722 430
rect 94838 400 95730 430
rect 95846 400 97074 430
rect 97190 400 98082 430
rect 98198 400 99426 430
rect 99542 400 100770 430
rect 100886 400 101778 430
rect 101894 400 103122 430
rect 103238 400 104466 430
rect 104582 400 105474 430
rect 105590 400 106818 430
rect 106934 400 107826 430
rect 107942 400 109170 430
rect 109286 400 110514 430
rect 110630 400 111522 430
rect 111638 400 112866 430
rect 112982 400 113874 430
rect 113990 400 115218 430
rect 115334 400 116562 430
rect 116678 400 117570 430
rect 117686 400 118914 430
rect 119030 400 120258 430
rect 120374 400 121266 430
rect 121382 400 122610 430
rect 122726 400 123578 430
<< metal3 >>
rect 100 124992 400 125048
rect 123800 124656 124100 124712
rect 100 123648 400 123704
rect 123800 123312 124100 123368
rect 100 122640 400 122696
rect 123800 122304 124100 122360
rect 100 121296 400 121352
rect 123800 120960 124100 121016
rect 100 120288 400 120344
rect 123800 119616 124100 119672
rect 100 118944 400 119000
rect 123800 118608 124100 118664
rect 100 117600 400 117656
rect 123800 117264 124100 117320
rect 100 116592 400 116648
rect 123800 116256 124100 116312
rect 100 115248 400 115304
rect 123800 114912 124100 114968
rect 100 113904 400 113960
rect 123800 113568 124100 113624
rect 100 112896 400 112952
rect 123800 112560 124100 112616
rect 100 111552 400 111608
rect 123800 111216 124100 111272
rect 100 110544 400 110600
rect 123800 109872 124100 109928
rect 100 109200 400 109256
rect 123800 108864 124100 108920
rect 100 107856 400 107912
rect 123800 107520 124100 107576
rect 100 106848 400 106904
rect 123800 106512 124100 106568
rect 100 105504 400 105560
rect 123800 105168 124100 105224
rect 100 104496 400 104552
rect 123800 103824 124100 103880
rect 100 103152 400 103208
rect 123800 102816 124100 102872
rect 100 101808 400 101864
rect 123800 101472 124100 101528
rect 100 100800 400 100856
rect 123800 100464 124100 100520
rect 100 99456 400 99512
rect 123800 99120 124100 99176
rect 100 98112 400 98168
rect 123800 97776 124100 97832
rect 100 97104 400 97160
rect 123800 96768 124100 96824
rect 100 95760 400 95816
rect 123800 95424 124100 95480
rect 100 94752 400 94808
rect 123800 94080 124100 94136
rect 100 93408 400 93464
rect 123800 93072 124100 93128
rect 100 92064 400 92120
rect 123800 91728 124100 91784
rect 100 91056 400 91112
rect 123800 90720 124100 90776
rect 100 89712 400 89768
rect 123800 89376 124100 89432
rect 100 88704 400 88760
rect 123800 88032 124100 88088
rect 100 87360 400 87416
rect 123800 87024 124100 87080
rect 100 86016 400 86072
rect 123800 85680 124100 85736
rect 100 85008 400 85064
rect 123800 84672 124100 84728
rect 100 83664 400 83720
rect 123800 83328 124100 83384
rect 100 82320 400 82376
rect 123800 81984 124100 82040
rect 100 81312 400 81368
rect 123800 80976 124100 81032
rect 100 79968 400 80024
rect 123800 79632 124100 79688
rect 100 78960 400 79016
rect 123800 78288 124100 78344
rect 100 77616 400 77672
rect 123800 77280 124100 77336
rect 100 76272 400 76328
rect 123800 75936 124100 75992
rect 100 75264 400 75320
rect 123800 74928 124100 74984
rect 100 73920 400 73976
rect 123800 73584 124100 73640
rect 100 72576 400 72632
rect 123800 72240 124100 72296
rect 100 71568 400 71624
rect 123800 71232 124100 71288
rect 100 70224 400 70280
rect 123800 69888 124100 69944
rect 100 69216 400 69272
rect 123800 68880 124100 68936
rect 100 67872 400 67928
rect 123800 67536 124100 67592
rect 100 66528 400 66584
rect 123800 66192 124100 66248
rect 100 65520 400 65576
rect 123800 65184 124100 65240
rect 100 64176 400 64232
rect 123800 63840 124100 63896
rect 100 63168 400 63224
rect 123800 62496 124100 62552
rect 100 61824 400 61880
rect 123800 61488 124100 61544
rect 100 60480 400 60536
rect 123800 60144 124100 60200
rect 100 59472 400 59528
rect 123800 59136 124100 59192
rect 100 58128 400 58184
rect 123800 57792 124100 57848
rect 100 56784 400 56840
rect 123800 56448 124100 56504
rect 100 55776 400 55832
rect 123800 55440 124100 55496
rect 100 54432 400 54488
rect 123800 54096 124100 54152
rect 100 53424 400 53480
rect 123800 53088 124100 53144
rect 100 52080 400 52136
rect 123800 51744 124100 51800
rect 100 50736 400 50792
rect 123800 50400 124100 50456
rect 100 49728 400 49784
rect 123800 49392 124100 49448
rect 100 48384 400 48440
rect 123800 48048 124100 48104
rect 100 47376 400 47432
rect 123800 46704 124100 46760
rect 100 46032 400 46088
rect 123800 45696 124100 45752
rect 100 44688 400 44744
rect 123800 44352 124100 44408
rect 100 43680 400 43736
rect 123800 43344 124100 43400
rect 100 42336 400 42392
rect 123800 42000 124100 42056
rect 100 40992 400 41048
rect 123800 40656 124100 40712
rect 100 39984 400 40040
rect 123800 39648 124100 39704
rect 100 38640 400 38696
rect 123800 38304 124100 38360
rect 100 37632 400 37688
rect 123800 36960 124100 37016
rect 100 36288 400 36344
rect 123800 35952 124100 36008
rect 100 34944 400 35000
rect 123800 34608 124100 34664
rect 100 33936 400 33992
rect 123800 33600 124100 33656
rect 100 32592 400 32648
rect 123800 32256 124100 32312
rect 100 31584 400 31640
rect 123800 30912 124100 30968
rect 100 30240 400 30296
rect 123800 29904 124100 29960
rect 100 28896 400 28952
rect 123800 28560 124100 28616
rect 100 27888 400 27944
rect 123800 27552 124100 27608
rect 100 26544 400 26600
rect 123800 26208 124100 26264
rect 100 25200 400 25256
rect 123800 24864 124100 24920
rect 100 24192 400 24248
rect 123800 23856 124100 23912
rect 100 22848 400 22904
rect 123800 22512 124100 22568
rect 100 21840 400 21896
rect 123800 21168 124100 21224
rect 100 20496 400 20552
rect 123800 20160 124100 20216
rect 100 19152 400 19208
rect 123800 18816 124100 18872
rect 100 18144 400 18200
rect 123800 17808 124100 17864
rect 100 16800 400 16856
rect 123800 16464 124100 16520
rect 100 15792 400 15848
rect 123800 15120 124100 15176
rect 100 14448 400 14504
rect 123800 14112 124100 14168
rect 100 13104 400 13160
rect 123800 12768 124100 12824
rect 100 12096 400 12152
rect 123800 11760 124100 11816
rect 100 10752 400 10808
rect 123800 10416 124100 10472
rect 100 9408 400 9464
rect 123800 9072 124100 9128
rect 100 8400 400 8456
rect 123800 8064 124100 8120
rect 100 7056 400 7112
rect 123800 6720 124100 6776
rect 100 6048 400 6104
rect 123800 5376 124100 5432
rect 100 4704 400 4760
rect 123800 4368 124100 4424
rect 100 3360 400 3416
rect 123800 3024 124100 3080
rect 100 2352 400 2408
rect 123800 2016 124100 2072
rect 100 1008 400 1064
rect 123800 672 124100 728
<< obsm3 >>
rect 9 123734 124194 124474
rect 9 123618 70 123734
rect 430 123618 124194 123734
rect 9 123398 124194 123618
rect 9 123282 123770 123398
rect 124130 123282 124194 123398
rect 9 122726 124194 123282
rect 9 122610 70 122726
rect 430 122610 124194 122726
rect 9 122390 124194 122610
rect 9 122274 123770 122390
rect 124130 122274 124194 122390
rect 9 121382 124194 122274
rect 9 121266 70 121382
rect 430 121266 124194 121382
rect 9 121046 124194 121266
rect 9 120930 123770 121046
rect 124130 120930 124194 121046
rect 9 120374 124194 120930
rect 9 120258 70 120374
rect 430 120258 124194 120374
rect 9 119702 124194 120258
rect 9 119586 123770 119702
rect 124130 119586 124194 119702
rect 9 119030 124194 119586
rect 9 118914 70 119030
rect 430 118914 124194 119030
rect 9 118694 124194 118914
rect 9 118578 123770 118694
rect 124130 118578 124194 118694
rect 9 117686 124194 118578
rect 9 117570 70 117686
rect 430 117570 124194 117686
rect 9 117350 124194 117570
rect 9 117234 123770 117350
rect 124130 117234 124194 117350
rect 9 116678 124194 117234
rect 9 116562 70 116678
rect 430 116562 124194 116678
rect 9 116342 124194 116562
rect 9 116226 123770 116342
rect 124130 116226 124194 116342
rect 9 115334 124194 116226
rect 9 115218 70 115334
rect 430 115218 124194 115334
rect 9 114998 124194 115218
rect 9 114882 123770 114998
rect 124130 114882 124194 114998
rect 9 113990 124194 114882
rect 9 113874 70 113990
rect 430 113874 124194 113990
rect 9 113654 124194 113874
rect 9 113538 123770 113654
rect 124130 113538 124194 113654
rect 9 112982 124194 113538
rect 9 112866 70 112982
rect 430 112866 124194 112982
rect 9 112646 124194 112866
rect 9 112530 123770 112646
rect 124130 112530 124194 112646
rect 9 111638 124194 112530
rect 9 111522 70 111638
rect 430 111522 124194 111638
rect 9 111302 124194 111522
rect 9 111186 123770 111302
rect 124130 111186 124194 111302
rect 9 110630 124194 111186
rect 9 110514 70 110630
rect 430 110514 124194 110630
rect 9 109958 124194 110514
rect 9 109842 123770 109958
rect 124130 109842 124194 109958
rect 9 109286 124194 109842
rect 9 109170 70 109286
rect 430 109170 124194 109286
rect 9 108950 124194 109170
rect 9 108834 123770 108950
rect 124130 108834 124194 108950
rect 9 107942 124194 108834
rect 9 107826 70 107942
rect 430 107826 124194 107942
rect 9 107606 124194 107826
rect 9 107490 123770 107606
rect 124130 107490 124194 107606
rect 9 106934 124194 107490
rect 9 106818 70 106934
rect 430 106818 124194 106934
rect 9 106598 124194 106818
rect 9 106482 123770 106598
rect 124130 106482 124194 106598
rect 9 105590 124194 106482
rect 9 105474 70 105590
rect 430 105474 124194 105590
rect 9 105254 124194 105474
rect 9 105138 123770 105254
rect 124130 105138 124194 105254
rect 9 104582 124194 105138
rect 9 104466 70 104582
rect 430 104466 124194 104582
rect 9 103910 124194 104466
rect 9 103794 123770 103910
rect 124130 103794 124194 103910
rect 9 103238 124194 103794
rect 9 103122 70 103238
rect 430 103122 124194 103238
rect 9 102902 124194 103122
rect 9 102786 123770 102902
rect 124130 102786 124194 102902
rect 9 101894 124194 102786
rect 9 101778 70 101894
rect 430 101778 124194 101894
rect 9 101558 124194 101778
rect 9 101442 123770 101558
rect 124130 101442 124194 101558
rect 9 100886 124194 101442
rect 9 100770 70 100886
rect 430 100770 124194 100886
rect 9 100550 124194 100770
rect 9 100434 123770 100550
rect 124130 100434 124194 100550
rect 9 99542 124194 100434
rect 9 99426 70 99542
rect 430 99426 124194 99542
rect 9 99206 124194 99426
rect 9 99090 123770 99206
rect 124130 99090 124194 99206
rect 9 98198 124194 99090
rect 9 98082 70 98198
rect 430 98082 124194 98198
rect 9 97862 124194 98082
rect 9 97746 123770 97862
rect 124130 97746 124194 97862
rect 9 97190 124194 97746
rect 9 97074 70 97190
rect 430 97074 124194 97190
rect 9 96854 124194 97074
rect 9 96738 123770 96854
rect 124130 96738 124194 96854
rect 9 95846 124194 96738
rect 9 95730 70 95846
rect 430 95730 124194 95846
rect 9 95510 124194 95730
rect 9 95394 123770 95510
rect 124130 95394 124194 95510
rect 9 94838 124194 95394
rect 9 94722 70 94838
rect 430 94722 124194 94838
rect 9 94166 124194 94722
rect 9 94050 123770 94166
rect 124130 94050 124194 94166
rect 9 93494 124194 94050
rect 9 93378 70 93494
rect 430 93378 124194 93494
rect 9 93158 124194 93378
rect 9 93042 123770 93158
rect 124130 93042 124194 93158
rect 9 92150 124194 93042
rect 9 92034 70 92150
rect 430 92034 124194 92150
rect 9 91814 124194 92034
rect 9 91698 123770 91814
rect 124130 91698 124194 91814
rect 9 91142 124194 91698
rect 9 91026 70 91142
rect 430 91026 124194 91142
rect 9 90806 124194 91026
rect 9 90690 123770 90806
rect 124130 90690 124194 90806
rect 9 89798 124194 90690
rect 9 89682 70 89798
rect 430 89682 124194 89798
rect 9 89462 124194 89682
rect 9 89346 123770 89462
rect 124130 89346 124194 89462
rect 9 88790 124194 89346
rect 9 88674 70 88790
rect 430 88674 124194 88790
rect 9 88118 124194 88674
rect 9 88002 123770 88118
rect 124130 88002 124194 88118
rect 9 87446 124194 88002
rect 9 87330 70 87446
rect 430 87330 124194 87446
rect 9 87110 124194 87330
rect 9 86994 123770 87110
rect 124130 86994 124194 87110
rect 9 86102 124194 86994
rect 9 85986 70 86102
rect 430 85986 124194 86102
rect 9 85766 124194 85986
rect 9 85650 123770 85766
rect 124130 85650 124194 85766
rect 9 85094 124194 85650
rect 9 84978 70 85094
rect 430 84978 124194 85094
rect 9 84758 124194 84978
rect 9 84642 123770 84758
rect 124130 84642 124194 84758
rect 9 83750 124194 84642
rect 9 83634 70 83750
rect 430 83634 124194 83750
rect 9 83414 124194 83634
rect 9 83298 123770 83414
rect 124130 83298 124194 83414
rect 9 82406 124194 83298
rect 9 82290 70 82406
rect 430 82290 124194 82406
rect 9 82070 124194 82290
rect 9 81954 123770 82070
rect 124130 81954 124194 82070
rect 9 81398 124194 81954
rect 9 81282 70 81398
rect 430 81282 124194 81398
rect 9 81062 124194 81282
rect 9 80946 123770 81062
rect 124130 80946 124194 81062
rect 9 80054 124194 80946
rect 9 79938 70 80054
rect 430 79938 124194 80054
rect 9 79718 124194 79938
rect 9 79602 123770 79718
rect 124130 79602 124194 79718
rect 9 79046 124194 79602
rect 9 78930 70 79046
rect 430 78930 124194 79046
rect 9 78374 124194 78930
rect 9 78258 123770 78374
rect 124130 78258 124194 78374
rect 9 77702 124194 78258
rect 9 77586 70 77702
rect 430 77586 124194 77702
rect 9 77366 124194 77586
rect 9 77250 123770 77366
rect 124130 77250 124194 77366
rect 9 76358 124194 77250
rect 9 76242 70 76358
rect 430 76242 124194 76358
rect 9 76022 124194 76242
rect 9 75906 123770 76022
rect 124130 75906 124194 76022
rect 9 75350 124194 75906
rect 9 75234 70 75350
rect 430 75234 124194 75350
rect 9 75014 124194 75234
rect 9 74898 123770 75014
rect 124130 74898 124194 75014
rect 9 74006 124194 74898
rect 9 73890 70 74006
rect 430 73890 124194 74006
rect 9 73670 124194 73890
rect 9 73554 123770 73670
rect 124130 73554 124194 73670
rect 9 72662 124194 73554
rect 9 72546 70 72662
rect 430 72546 124194 72662
rect 9 72326 124194 72546
rect 9 72210 123770 72326
rect 124130 72210 124194 72326
rect 9 71654 124194 72210
rect 9 71538 70 71654
rect 430 71538 124194 71654
rect 9 71318 124194 71538
rect 9 71202 123770 71318
rect 124130 71202 124194 71318
rect 9 70310 124194 71202
rect 9 70194 70 70310
rect 430 70194 124194 70310
rect 9 69974 124194 70194
rect 9 69858 123770 69974
rect 124130 69858 124194 69974
rect 9 69302 124194 69858
rect 9 69186 70 69302
rect 430 69186 124194 69302
rect 9 68966 124194 69186
rect 9 68850 123770 68966
rect 124130 68850 124194 68966
rect 9 67958 124194 68850
rect 9 67842 70 67958
rect 430 67842 124194 67958
rect 9 67622 124194 67842
rect 9 67506 123770 67622
rect 124130 67506 124194 67622
rect 9 66614 124194 67506
rect 9 66498 70 66614
rect 430 66498 124194 66614
rect 9 66278 124194 66498
rect 9 66162 123770 66278
rect 124130 66162 124194 66278
rect 9 65606 124194 66162
rect 9 65490 70 65606
rect 430 65490 124194 65606
rect 9 65270 124194 65490
rect 9 65154 123770 65270
rect 124130 65154 124194 65270
rect 9 64262 124194 65154
rect 9 64146 70 64262
rect 430 64146 124194 64262
rect 9 63926 124194 64146
rect 9 63810 123770 63926
rect 124130 63810 124194 63926
rect 9 63254 124194 63810
rect 9 63138 70 63254
rect 430 63138 124194 63254
rect 9 62582 124194 63138
rect 9 62466 123770 62582
rect 124130 62466 124194 62582
rect 9 61910 124194 62466
rect 9 61794 70 61910
rect 430 61794 124194 61910
rect 9 61574 124194 61794
rect 9 61458 123770 61574
rect 124130 61458 124194 61574
rect 9 60566 124194 61458
rect 9 60450 70 60566
rect 430 60450 124194 60566
rect 9 60230 124194 60450
rect 9 60114 123770 60230
rect 124130 60114 124194 60230
rect 9 59558 124194 60114
rect 9 59442 70 59558
rect 430 59442 124194 59558
rect 9 59222 124194 59442
rect 9 59106 123770 59222
rect 124130 59106 124194 59222
rect 9 58214 124194 59106
rect 9 58098 70 58214
rect 430 58098 124194 58214
rect 9 57878 124194 58098
rect 9 57762 123770 57878
rect 124130 57762 124194 57878
rect 9 56870 124194 57762
rect 9 56754 70 56870
rect 430 56754 124194 56870
rect 9 56534 124194 56754
rect 9 56418 123770 56534
rect 124130 56418 124194 56534
rect 9 55862 124194 56418
rect 9 55746 70 55862
rect 430 55746 124194 55862
rect 9 55526 124194 55746
rect 9 55410 123770 55526
rect 124130 55410 124194 55526
rect 9 54518 124194 55410
rect 9 54402 70 54518
rect 430 54402 124194 54518
rect 9 54182 124194 54402
rect 9 54066 123770 54182
rect 124130 54066 124194 54182
rect 9 53510 124194 54066
rect 9 53394 70 53510
rect 430 53394 124194 53510
rect 9 53174 124194 53394
rect 9 53058 123770 53174
rect 124130 53058 124194 53174
rect 9 52166 124194 53058
rect 9 52050 70 52166
rect 430 52050 124194 52166
rect 9 51830 124194 52050
rect 9 51714 123770 51830
rect 124130 51714 124194 51830
rect 9 50822 124194 51714
rect 9 50706 70 50822
rect 430 50706 124194 50822
rect 9 50486 124194 50706
rect 9 50370 123770 50486
rect 124130 50370 124194 50486
rect 9 49814 124194 50370
rect 9 49698 70 49814
rect 430 49698 124194 49814
rect 9 49478 124194 49698
rect 9 49362 123770 49478
rect 124130 49362 124194 49478
rect 9 48470 124194 49362
rect 9 48354 70 48470
rect 430 48354 124194 48470
rect 9 48134 124194 48354
rect 9 48018 123770 48134
rect 124130 48018 124194 48134
rect 9 47462 124194 48018
rect 9 47346 70 47462
rect 430 47346 124194 47462
rect 9 46790 124194 47346
rect 9 46674 123770 46790
rect 124130 46674 124194 46790
rect 9 46118 124194 46674
rect 9 46002 70 46118
rect 430 46002 124194 46118
rect 9 45782 124194 46002
rect 9 45666 123770 45782
rect 124130 45666 124194 45782
rect 9 44774 124194 45666
rect 9 44658 70 44774
rect 430 44658 124194 44774
rect 9 44438 124194 44658
rect 9 44322 123770 44438
rect 124130 44322 124194 44438
rect 9 43766 124194 44322
rect 9 43650 70 43766
rect 430 43650 124194 43766
rect 9 43430 124194 43650
rect 9 43314 123770 43430
rect 124130 43314 124194 43430
rect 9 42422 124194 43314
rect 9 42306 70 42422
rect 430 42306 124194 42422
rect 9 42086 124194 42306
rect 9 41970 123770 42086
rect 124130 41970 124194 42086
rect 9 41078 124194 41970
rect 9 40962 70 41078
rect 430 40962 124194 41078
rect 9 40742 124194 40962
rect 9 40626 123770 40742
rect 124130 40626 124194 40742
rect 9 40070 124194 40626
rect 9 39954 70 40070
rect 430 39954 124194 40070
rect 9 39734 124194 39954
rect 9 39618 123770 39734
rect 124130 39618 124194 39734
rect 9 38726 124194 39618
rect 9 38610 70 38726
rect 430 38610 124194 38726
rect 9 38390 124194 38610
rect 9 38274 123770 38390
rect 124130 38274 124194 38390
rect 9 37718 124194 38274
rect 9 37602 70 37718
rect 430 37602 124194 37718
rect 9 37046 124194 37602
rect 9 36930 123770 37046
rect 124130 36930 124194 37046
rect 9 36374 124194 36930
rect 9 36258 70 36374
rect 430 36258 124194 36374
rect 9 36038 124194 36258
rect 9 35922 123770 36038
rect 124130 35922 124194 36038
rect 9 35030 124194 35922
rect 9 34914 70 35030
rect 430 34914 124194 35030
rect 9 34694 124194 34914
rect 9 34578 123770 34694
rect 124130 34578 124194 34694
rect 9 34022 124194 34578
rect 9 33906 70 34022
rect 430 33906 124194 34022
rect 9 33686 124194 33906
rect 9 33570 123770 33686
rect 124130 33570 124194 33686
rect 9 32678 124194 33570
rect 9 32562 70 32678
rect 430 32562 124194 32678
rect 9 32342 124194 32562
rect 9 32226 123770 32342
rect 124130 32226 124194 32342
rect 9 31670 124194 32226
rect 9 31554 70 31670
rect 430 31554 124194 31670
rect 9 30998 124194 31554
rect 9 30882 123770 30998
rect 124130 30882 124194 30998
rect 9 30326 124194 30882
rect 9 30210 70 30326
rect 430 30210 124194 30326
rect 9 29990 124194 30210
rect 9 29874 123770 29990
rect 124130 29874 124194 29990
rect 9 28982 124194 29874
rect 9 28866 70 28982
rect 430 28866 124194 28982
rect 9 28646 124194 28866
rect 9 28530 123770 28646
rect 124130 28530 124194 28646
rect 9 27974 124194 28530
rect 9 27858 70 27974
rect 430 27858 124194 27974
rect 9 27638 124194 27858
rect 9 27522 123770 27638
rect 124130 27522 124194 27638
rect 9 26630 124194 27522
rect 9 26514 70 26630
rect 430 26514 124194 26630
rect 9 26294 124194 26514
rect 9 26178 123770 26294
rect 124130 26178 124194 26294
rect 9 25286 124194 26178
rect 9 25170 70 25286
rect 430 25170 124194 25286
rect 9 24950 124194 25170
rect 9 24834 123770 24950
rect 124130 24834 124194 24950
rect 9 24278 124194 24834
rect 9 24162 70 24278
rect 430 24162 124194 24278
rect 9 23942 124194 24162
rect 9 23826 123770 23942
rect 124130 23826 124194 23942
rect 9 22934 124194 23826
rect 9 22818 70 22934
rect 430 22818 124194 22934
rect 9 22598 124194 22818
rect 9 22482 123770 22598
rect 124130 22482 124194 22598
rect 9 21926 124194 22482
rect 9 21810 70 21926
rect 430 21810 124194 21926
rect 9 21254 124194 21810
rect 9 21138 123770 21254
rect 124130 21138 124194 21254
rect 9 20582 124194 21138
rect 9 20466 70 20582
rect 430 20466 124194 20582
rect 9 20246 124194 20466
rect 9 20130 123770 20246
rect 124130 20130 124194 20246
rect 9 19238 124194 20130
rect 9 19122 70 19238
rect 430 19122 124194 19238
rect 9 18902 124194 19122
rect 9 18786 123770 18902
rect 124130 18786 124194 18902
rect 9 18230 124194 18786
rect 9 18114 70 18230
rect 430 18114 124194 18230
rect 9 17894 124194 18114
rect 9 17778 123770 17894
rect 124130 17778 124194 17894
rect 9 16886 124194 17778
rect 9 16770 70 16886
rect 430 16770 124194 16886
rect 9 16550 124194 16770
rect 9 16434 123770 16550
rect 124130 16434 124194 16550
rect 9 15878 124194 16434
rect 9 15762 70 15878
rect 430 15762 124194 15878
rect 9 15206 124194 15762
rect 9 15090 123770 15206
rect 124130 15090 124194 15206
rect 9 14534 124194 15090
rect 9 14418 70 14534
rect 430 14418 124194 14534
rect 9 14198 124194 14418
rect 9 14082 123770 14198
rect 124130 14082 124194 14198
rect 9 13190 124194 14082
rect 9 13074 70 13190
rect 430 13074 124194 13190
rect 9 12854 124194 13074
rect 9 12738 123770 12854
rect 124130 12738 124194 12854
rect 9 12182 124194 12738
rect 9 12066 70 12182
rect 430 12066 124194 12182
rect 9 11846 124194 12066
rect 9 11730 123770 11846
rect 124130 11730 124194 11846
rect 9 10838 124194 11730
rect 9 10722 70 10838
rect 430 10722 124194 10838
rect 9 10502 124194 10722
rect 9 10386 123770 10502
rect 124130 10386 124194 10502
rect 9 9494 124194 10386
rect 9 9378 70 9494
rect 430 9378 124194 9494
rect 9 9158 124194 9378
rect 9 9042 123770 9158
rect 124130 9042 124194 9158
rect 9 8486 124194 9042
rect 9 8370 70 8486
rect 430 8370 124194 8486
rect 9 8150 124194 8370
rect 9 8034 123770 8150
rect 124130 8034 124194 8150
rect 9 7142 124194 8034
rect 9 7026 70 7142
rect 430 7026 124194 7142
rect 9 6806 124194 7026
rect 9 6690 123770 6806
rect 124130 6690 124194 6806
rect 9 6134 124194 6690
rect 9 6018 70 6134
rect 430 6018 124194 6134
rect 9 5462 124194 6018
rect 9 5346 123770 5462
rect 124130 5346 124194 5462
rect 9 4790 124194 5346
rect 9 4674 70 4790
rect 430 4674 124194 4790
rect 9 4454 124194 4674
rect 9 4338 123770 4454
rect 124130 4338 124194 4454
rect 9 3446 124194 4338
rect 9 3330 70 3446
rect 430 3330 124194 3446
rect 9 3110 124194 3330
rect 9 2994 123770 3110
rect 124130 2994 124194 3110
rect 9 2438 124194 2994
rect 9 2322 70 2438
rect 430 2322 124194 2438
rect 9 2102 124194 2322
rect 9 1986 123770 2102
rect 124130 1986 124194 2102
rect 9 1094 124194 1986
rect 9 978 70 1094
rect 430 978 124194 1094
rect 9 798 124194 978
<< metal4 >>
rect 2224 1538 2384 124294
rect 9904 1538 10064 124294
rect 17584 1538 17744 124294
rect 25264 1538 25424 124294
rect 32944 1538 33104 124294
rect 40624 1538 40784 124294
rect 48304 1538 48464 124294
rect 55984 1538 56144 124294
rect 63664 1538 63824 124294
rect 71344 1538 71504 124294
rect 79024 1538 79184 124294
rect 86704 1538 86864 124294
rect 94384 1538 94544 124294
rect 102064 1538 102224 124294
rect 109744 1538 109904 124294
rect 117424 1538 117584 124294
<< obsm4 >>
rect 2142 1508 2194 124087
rect 2414 1508 9874 124087
rect 10094 1508 17554 124087
rect 17774 1508 25234 124087
rect 25454 1508 32914 124087
rect 33134 1508 40594 124087
rect 40814 1508 48274 124087
rect 48494 1508 55954 124087
rect 56174 1508 63634 124087
rect 63854 1508 71314 124087
rect 71534 1508 78994 124087
rect 79214 1508 86674 124087
rect 86894 1508 94354 124087
rect 94574 1508 102034 124087
rect 102254 1508 109714 124087
rect 109934 1508 117394 124087
rect 117614 1508 122626 124087
rect 2142 1353 122626 1508
<< labels >>
rlabel metal2 s 73248 125592 73304 125892 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 16128 125592 16184 125892 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 94752 400 94808 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 123800 124656 124100 124712 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 8400 400 8456 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 91392 125592 91448 125892 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 123800 80976 124100 81032 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 100 58128 400 58184 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 123800 45696 124100 45752 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 100 124992 400 125048 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 121632 125592 121688 125892 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 100 99456 400 99512 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 123800 20160 124100 20216 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 100 64176 400 64232 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 26880 125592 26936 125892 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 100 111552 400 111608 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 106848 100 106904 400 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 123800 26208 124100 26264 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 121296 100 121352 400 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 6048 400 6104 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 122976 125592 123032 125892 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 63504 125592 63560 125892 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 100 13104 400 13160 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 100 24192 400 24248 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 59808 125592 59864 125892 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 123800 120960 124100 121016 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 13440 125592 13496 125892 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 123800 94080 124100 94136 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 100 71568 400 71624 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 105840 125592 105896 125892 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 123800 30912 124100 30968 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 123800 53088 124100 53144 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 10080 125592 10136 125892 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 101136 125592 101192 125892 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 43680 100 43736 400 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 123800 96768 124100 96824 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 25200 100 25256 400 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 123800 11760 124100 11816 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 123800 21168 124100 21224 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 92064 100 92120 400 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 68208 125592 68264 125892 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 121296 400 121352 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 100 2352 400 2408 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 20832 125592 20888 125892 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 32928 125592 32984 125892 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 17136 125592 17192 125892 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 93408 400 93464 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 73920 100 73976 400 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 123800 108864 124100 108920 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 123800 27552 124100 27608 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 100 95760 400 95816 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 116592 100 116648 400 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 100 107856 400 107912 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 103152 100 103208 400 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 53760 125592 53816 125892 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 67200 125592 67256 125892 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 111552 100 111608 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 123800 44352 124100 44408 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 90048 125592 90104 125892 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 104832 125592 104888 125892 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 12096 100 12152 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 117936 125592 117992 125892 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 49728 100 49784 400 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 18480 125592 18536 125892 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 5040 125592 5096 125892 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 100 55776 400 55832 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 104496 100 104552 400 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 123800 49392 124100 49448 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 109536 125592 109592 125892 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 42336 400 42392 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 123800 18816 124100 18872 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 114576 125592 114632 125892 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 52080 100 52136 400 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 77616 100 77672 400 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 123800 14112 124100 14168 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 123800 78288 124100 78344 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 100 85008 400 85064 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 123800 113568 124100 113624 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 56112 125592 56168 125892 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 14448 100 14504 400 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 83664 400 83720 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 79968 100 80024 400 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 8400 100 8456 400 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 123800 71232 124100 71288 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 55776 100 55832 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 40992 100 41048 400 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 123800 40656 124100 40712 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 105504 100 105560 400 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 50736 400 50792 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 116928 125592 116984 125892 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 123648 400 123704 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 100 65520 400 65576 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 82320 100 82376 400 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 70560 125592 70616 125892 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 100 78960 400 79016 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 123800 24864 124100 24920 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 100 56784 400 56840 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 81312 100 81368 400 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 123800 17808 124100 17864 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 123800 123312 124100 123368 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 123800 4368 124100 4424 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 28224 125592 28280 125892 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 60816 125592 60872 125892 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 100 52080 400 52136 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 72576 400 72632 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 76608 125592 76664 125892 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 89712 100 89768 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 11088 125592 11144 125892 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 37632 400 37688 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 122640 100 122696 400 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46032 100 46088 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 37632 100 37688 400 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 51408 125592 51464 125892 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 113232 125592 113288 125892 6 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 58128 100 58184 400 6 la_data_in[11]
port 117 nsew signal input
rlabel metal3 s 100 76272 400 76328 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 97440 125592 97496 125892 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 123800 122304 124100 122360 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 123800 32256 124100 32312 6 la_data_in[15]
port 121 nsew signal input
rlabel metal3 s 100 81312 400 81368 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 123800 23856 124100 23912 6 la_data_in[17]
port 123 nsew signal input
rlabel metal3 s 100 12096 400 12152 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 7056 400 7112 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 99792 125592 99848 125892 6 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 77952 125592 78008 125892 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 123800 103824 124100 103880 6 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 92400 125592 92456 125892 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 100 36288 400 36344 6 la_data_in[23]
port 130 nsew signal input
rlabel metal3 s 100 60480 400 60536 6 la_data_in[24]
port 131 nsew signal input
rlabel metal3 s 100 106848 400 106904 6 la_data_in[25]
port 132 nsew signal input
rlabel metal3 s 123800 114912 124100 114968 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 123800 68880 124100 68936 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 122640 400 122696 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 123800 51744 124100 51800 6 la_data_in[29]
port 136 nsew signal input
rlabel metal3 s 123800 107520 124100 107576 6 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 117600 100 117656 400 6 la_data_in[30]
port 138 nsew signal input
rlabel metal3 s 100 28896 400 28952 6 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 87360 100 87416 400 6 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 45024 125592 45080 125892 6 la_data_in[33]
port 141 nsew signal input
rlabel metal3 s 100 86016 400 86072 6 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 52416 125592 52472 125892 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 84000 125592 84056 125892 6 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 42336 100 42392 400 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 59472 100 59528 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal3 s 100 118944 400 119000 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 100 53424 400 53480 6 la_data_in[3]
port 148 nsew signal input
rlabel metal3 s 100 88704 400 88760 6 la_data_in[40]
port 149 nsew signal input
rlabel metal3 s 123800 90720 124100 90776 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 123800 89376 124100 89432 6 la_data_in[42]
port 151 nsew signal input
rlabel metal3 s 100 10752 400 10808 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 100 32592 400 32648 6 la_data_in[44]
port 153 nsew signal input
rlabel metal3 s 100 9408 400 9464 6 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 30240 100 30296 400 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 50064 125592 50120 125892 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 56784 100 56840 400 6 la_data_in[48]
port 157 nsew signal input
rlabel metal3 s 100 113904 400 113960 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 37968 125592 38024 125892 6 la_data_in[4]
port 159 nsew signal input
rlabel metal3 s 123800 33600 124100 33656 6 la_data_in[50]
port 160 nsew signal input
rlabel metal3 s 100 33936 400 33992 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 100 34944 400 35000 6 la_data_in[52]
port 162 nsew signal input
rlabel metal3 s 123800 3024 124100 3080 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 44688 100 44744 400 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 48384 400 48440 6 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 21840 100 21896 400 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 86352 125592 86408 125892 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 95088 125592 95144 125892 6 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 72576 100 72632 400 6 la_data_in[59]
port 169 nsew signal input
rlabel metal3 s 123800 60144 124100 60200 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 100 61824 400 61880 6 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 336 125592 392 125892 6 la_data_in[61]
port 172 nsew signal input
rlabel metal3 s 100 104496 400 104552 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 69552 125592 69608 125892 6 la_data_in[63]
port 174 nsew signal input
rlabel metal3 s 100 18144 400 18200 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 100 77616 400 77672 6 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 88704 100 88760 400 6 la_data_in[8]
port 177 nsew signal input
rlabel metal3 s 100 91056 400 91112 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 35280 125592 35336 125892 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 123800 50400 124100 50456 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 123800 117264 124100 117320 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 123800 67536 124100 67592 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 62160 125592 62216 125892 6 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 54768 125592 54824 125892 6 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 65520 100 65576 400 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 123800 57792 124100 57848 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 58464 125592 58520 125892 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 123800 87024 124100 87080 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 65856 125592 65912 125892 6 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 36288 100 36344 400 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 100 19152 400 19208 6 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 66528 100 66584 400 6 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 108192 125592 108248 125892 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 16800 100 16856 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 16800 400 16856 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 53424 100 53480 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 98112 400 98168 6 la_data_out[26]
port 197 nsew signal output
rlabel metal3 s 123800 56448 124100 56504 6 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 3696 125592 3752 125892 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 19488 125592 19544 125892 6 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 2688 125592 2744 125892 6 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 60480 100 60536 400 6 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 33936 100 33992 400 6 la_data_out[31]
port 203 nsew signal output
rlabel metal3 s 123800 100464 124100 100520 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 123800 48048 124100 48104 6 la_data_out[33]
port 205 nsew signal output
rlabel metal3 s 123800 2016 124100 2072 6 la_data_out[34]
port 206 nsew signal output
rlabel metal3 s 123800 16464 124100 16520 6 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 87696 125592 87752 125892 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 100 112896 400 112952 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 123800 36960 124100 37016 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 123800 105168 124100 105224 6 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 7056 100 7112 400 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 50736 100 50792 400 6 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 75600 125592 75656 125892 6 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 113904 100 113960 400 6 la_data_out[42]
port 215 nsew signal output
rlabel metal3 s 100 89712 400 89768 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 28896 100 28952 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 112896 100 112952 400 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 71904 125592 71960 125892 6 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 44016 125592 44072 125892 6 la_data_out[47]
port 220 nsew signal output
rlabel metal3 s 100 46032 400 46088 6 la_data_out[48]
port 221 nsew signal output
rlabel metal3 s 123800 8064 124100 8120 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 69216 100 69272 400 6 la_data_out[4]
port 223 nsew signal output
rlabel metal3 s 100 117600 400 117656 6 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 47712 125592 47768 125892 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 123800 28560 124100 28616 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 100800 400 100856 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 123800 85680 124100 85736 6 la_data_out[54]
port 228 nsew signal output
rlabel metal3 s 123800 111216 124100 111272 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 123800 74928 124100 74984 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 102144 125592 102200 125892 6 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 32592 100 32648 400 6 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 107856 100 107912 400 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 123800 9072 124100 9128 6 la_data_out[5]
port 234 nsew signal output
rlabel metal3 s 100 87360 400 87416 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 120624 125592 120680 125892 6 la_data_out[61]
port 236 nsew signal output
rlabel metal3 s 100 116592 400 116648 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 123800 59136 124100 59192 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 123800 46704 124100 46760 6 la_data_out[6]
port 239 nsew signal output
rlabel metal3 s 123800 88032 124100 88088 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 123800 69888 124100 69944 6 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 48720 125592 48776 125892 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 100 44688 400 44744 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 100 4704 400 4760 6 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 109200 100 109256 400 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 18144 100 18200 400 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 15792 400 15848 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 8736 125592 8792 125892 6 la_oenb[14]
port 248 nsew signal input
rlabel metal3 s 123800 10416 124100 10472 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 24528 125592 24584 125892 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 110544 400 110600 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 22176 125592 22232 125892 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 100 3360 400 3416 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 34944 100 35000 400 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 31584 400 31640 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 110544 100 110600 400 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 25872 125592 25928 125892 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 22848 100 22904 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 123800 65184 124100 65240 6 la_oenb[24]
port 259 nsew signal input
rlabel metal3 s 123800 118608 124100 118664 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 123984 125592 124040 125892 6 la_oenb[26]
port 261 nsew signal input
rlabel metal3 s 123800 106512 124100 106568 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 123800 102816 124100 102872 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 123800 101472 124100 101528 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 63168 100 63224 400 6 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 111888 125592 111944 125892 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 3360 100 3416 400 6 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 1008 100 1064 400 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 1344 125592 1400 125892 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 64176 100 64232 400 6 la_oenb[34]
port 270 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 la_oenb[35]
port 271 nsew signal input
rlabel metal3 s 100 69216 400 69272 6 la_oenb[36]
port 272 nsew signal input
rlabel metal3 s 100 39984 400 40040 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 46368 125592 46424 125892 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 79968 400 80024 6 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 24192 100 24248 400 6 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 54432 100 54488 400 6 la_oenb[40]
port 277 nsew signal input
rlabel metal3 s 100 63168 400 63224 6 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 99456 100 99512 400 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 47376 100 47432 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal3 s 100 92064 400 92120 6 la_oenb[44]
port 281 nsew signal input
rlabel metal3 s 123800 61488 124100 61544 6 la_oenb[45]
port 282 nsew signal input
rlabel metal3 s 123800 83328 124100 83384 6 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 95760 100 95816 400 6 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 40320 125592 40376 125892 6 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 123648 100 123704 400 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 123800 79632 124100 79688 6 la_oenb[4]
port 287 nsew signal input
rlabel metal3 s 100 75264 400 75320 6 la_oenb[50]
port 288 nsew signal input
rlabel metal3 s 123800 63840 124100 63896 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 94752 100 94808 400 6 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 110880 125592 110936 125892 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 123800 12768 124100 12824 6 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 74256 125592 74312 125892 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 115248 100 115304 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 30576 125592 30632 125892 6 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 15792 100 15848 400 6 la_oenb[58]
port 296 nsew signal input
rlabel metal3 s 100 1008 400 1064 6 la_oenb[59]
port 297 nsew signal input
rlabel metal3 s 100 120288 400 120344 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 123800 81984 124100 82040 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 31584 100 31640 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 118944 100 119000 400 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 22848 400 22904 6 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 107184 125592 107240 125892 6 la_oenb[6]
port 303 nsew signal input
rlabel metal3 s 123800 95424 124100 95480 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 31920 125592 31976 125892 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 42672 125592 42728 125892 6 la_oenb[9]
port 306 nsew signal input
rlabel metal4 s 2224 1538 2384 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 124294 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 124294 6 vss
port 308 nsew ground bidirectional
rlabel metal3 s 123800 22512 124100 22568 6 wb_clk_i
port 309 nsew signal input
rlabel metal2 s 23184 125592 23240 125892 6 wb_rst_i
port 310 nsew signal input
rlabel metal3 s 123800 43344 124100 43400 6 wbs_ack_o
port 311 nsew signal output
rlabel metal2 s 82992 125592 83048 125892 6 wbs_adr_i[0]
port 312 nsew signal input
rlabel metal2 s 57456 125592 57512 125892 6 wbs_adr_i[10]
port 313 nsew signal input
rlabel metal2 s 7392 125592 7448 125892 6 wbs_adr_i[11]
port 314 nsew signal input
rlabel metal2 s 10752 100 10808 400 6 wbs_adr_i[12]
port 315 nsew signal input
rlabel metal3 s 100 30240 400 30296 6 wbs_adr_i[13]
port 316 nsew signal input
rlabel metal3 s 123800 91728 124100 91784 6 wbs_adr_i[14]
port 317 nsew signal input
rlabel metal3 s 123800 84672 124100 84728 6 wbs_adr_i[15]
port 318 nsew signal input
rlabel metal2 s 78960 100 79016 400 6 wbs_adr_i[16]
port 319 nsew signal input
rlabel metal3 s 100 70224 400 70280 6 wbs_adr_i[17]
port 320 nsew signal input
rlabel metal3 s 123800 39648 124100 39704 6 wbs_adr_i[18]
port 321 nsew signal input
rlabel metal2 s 120288 100 120344 400 6 wbs_adr_i[19]
port 322 nsew signal input
rlabel metal2 s 80304 125592 80360 125892 6 wbs_adr_i[1]
port 323 nsew signal input
rlabel metal3 s 100 67872 400 67928 6 wbs_adr_i[20]
port 324 nsew signal input
rlabel metal2 s 70224 100 70280 400 6 wbs_adr_i[21]
port 325 nsew signal input
rlabel metal2 s 100800 100 100856 400 6 wbs_adr_i[22]
port 326 nsew signal input
rlabel metal3 s 123800 29904 124100 29960 6 wbs_adr_i[23]
port 327 nsew signal input
rlabel metal2 s 14784 125592 14840 125892 6 wbs_adr_i[24]
port 328 nsew signal input
rlabel metal3 s 100 21840 400 21896 6 wbs_adr_i[25]
port 329 nsew signal input
rlabel metal2 s 13104 100 13160 400 6 wbs_adr_i[26]
port 330 nsew signal input
rlabel metal2 s 41664 125592 41720 125892 6 wbs_adr_i[27]
port 331 nsew signal input
rlabel metal3 s 123800 73584 124100 73640 6 wbs_adr_i[28]
port 332 nsew signal input
rlabel metal3 s 123800 119616 124100 119672 6 wbs_adr_i[29]
port 333 nsew signal input
rlabel metal3 s 100 14448 400 14504 6 wbs_adr_i[2]
port 334 nsew signal input
rlabel metal3 s 100 49728 400 49784 6 wbs_adr_i[30]
port 335 nsew signal input
rlabel metal3 s 123800 54096 124100 54152 6 wbs_adr_i[31]
port 336 nsew signal input
rlabel metal2 s 97104 100 97160 400 6 wbs_adr_i[3]
port 337 nsew signal input
rlabel metal2 s 96096 125592 96152 125892 6 wbs_adr_i[4]
port 338 nsew signal input
rlabel metal2 s 93408 100 93464 400 6 wbs_adr_i[5]
port 339 nsew signal input
rlabel metal2 s 39984 100 40040 400 6 wbs_adr_i[6]
port 340 nsew signal input
rlabel metal2 s 6048 100 6104 400 6 wbs_adr_i[7]
port 341 nsew signal input
rlabel metal3 s 123800 672 124100 728 6 wbs_adr_i[8]
port 342 nsew signal input
rlabel metal3 s 123800 34608 124100 34664 6 wbs_adr_i[9]
port 343 nsew signal input
rlabel metal2 s 38976 125592 39032 125892 6 wbs_cyc_i
port 344 nsew signal input
rlabel metal3 s 123800 109872 124100 109928 6 wbs_dat_i[0]
port 345 nsew signal input
rlabel metal3 s 100 97104 400 97160 6 wbs_dat_i[10]
port 346 nsew signal input
rlabel metal3 s 100 105504 400 105560 6 wbs_dat_i[11]
port 347 nsew signal input
rlabel metal3 s 100 101808 400 101864 6 wbs_dat_i[12]
port 348 nsew signal input
rlabel metal2 s 4704 100 4760 400 6 wbs_dat_i[13]
port 349 nsew signal input
rlabel metal3 s 100 26544 400 26600 6 wbs_dat_i[14]
port 350 nsew signal input
rlabel metal3 s 123800 66192 124100 66248 6 wbs_dat_i[15]
port 351 nsew signal input
rlabel metal2 s 71568 100 71624 400 6 wbs_dat_i[16]
port 352 nsew signal input
rlabel metal3 s 100 20496 400 20552 6 wbs_dat_i[17]
port 353 nsew signal input
rlabel metal2 s 115584 125592 115640 125892 6 wbs_dat_i[18]
port 354 nsew signal input
rlabel metal2 s 6384 125592 6440 125892 6 wbs_dat_i[19]
port 355 nsew signal input
rlabel metal2 s 19152 100 19208 400 6 wbs_dat_i[1]
port 356 nsew signal input
rlabel metal3 s 123800 75936 124100 75992 6 wbs_dat_i[20]
port 357 nsew signal input
rlabel metal2 s 119280 125592 119336 125892 6 wbs_dat_i[21]
port 358 nsew signal input
rlabel metal3 s 100 73920 400 73976 6 wbs_dat_i[22]
port 359 nsew signal input
rlabel metal3 s 123800 99120 124100 99176 6 wbs_dat_i[23]
port 360 nsew signal input
rlabel metal3 s 123800 42000 124100 42056 6 wbs_dat_i[24]
port 361 nsew signal input
rlabel metal2 s 86016 100 86072 400 6 wbs_dat_i[25]
port 362 nsew signal input
rlabel metal2 s 103488 125592 103544 125892 6 wbs_dat_i[26]
port 363 nsew signal input
rlabel metal2 s 29232 125592 29288 125892 6 wbs_dat_i[27]
port 364 nsew signal input
rlabel metal2 s 38640 100 38696 400 6 wbs_dat_i[28]
port 365 nsew signal input
rlabel metal3 s 123800 77280 124100 77336 6 wbs_dat_i[29]
port 366 nsew signal input
rlabel metal2 s 101808 100 101864 400 6 wbs_dat_i[2]
port 367 nsew signal input
rlabel metal3 s 123800 38304 124100 38360 6 wbs_dat_i[30]
port 368 nsew signal input
rlabel metal3 s 100 66528 400 66584 6 wbs_dat_i[31]
port 369 nsew signal input
rlabel metal3 s 123800 5376 124100 5432 6 wbs_dat_i[3]
port 370 nsew signal input
rlabel metal2 s 20496 100 20552 400 6 wbs_dat_i[4]
port 371 nsew signal input
rlabel metal2 s 61824 100 61880 400 6 wbs_dat_i[5]
port 372 nsew signal input
rlabel metal3 s 123800 55440 124100 55496 6 wbs_dat_i[6]
port 373 nsew signal input
rlabel metal2 s 98784 125592 98840 125892 6 wbs_dat_i[7]
port 374 nsew signal input
rlabel metal3 s 123800 112560 124100 112616 6 wbs_dat_i[8]
port 375 nsew signal input
rlabel metal3 s 123800 6720 124100 6776 6 wbs_dat_i[9]
port 376 nsew signal input
rlabel metal3 s 100 25200 400 25256 6 wbs_dat_o[0]
port 377 nsew signal output
rlabel metal3 s 123800 72240 124100 72296 6 wbs_dat_o[10]
port 378 nsew signal output
rlabel metal2 s 2352 100 2408 400 6 wbs_dat_o[11]
port 379 nsew signal output
rlabel metal3 s 123800 116256 124100 116312 6 wbs_dat_o[12]
port 380 nsew signal output
rlabel metal2 s 93744 125592 93800 125892 6 wbs_dat_o[13]
port 381 nsew signal output
rlabel metal3 s 123800 15120 124100 15176 6 wbs_dat_o[14]
port 382 nsew signal output
rlabel metal2 s 89040 125592 89096 125892 6 wbs_dat_o[15]
port 383 nsew signal output
rlabel metal2 s 85008 100 85064 400 6 wbs_dat_o[16]
port 384 nsew signal output
rlabel metal3 s 100 38640 400 38696 6 wbs_dat_o[17]
port 385 nsew signal output
rlabel metal2 s 83664 100 83720 400 6 wbs_dat_o[18]
port 386 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 387 nsew signal output
rlabel metal2 s 98112 100 98168 400 6 wbs_dat_o[1]
port 388 nsew signal output
rlabel metal3 s 100 59472 400 59528 6 wbs_dat_o[20]
port 389 nsew signal output
rlabel metal3 s 100 109200 400 109256 6 wbs_dat_o[21]
port 390 nsew signal output
rlabel metal2 s 34272 125592 34328 125892 6 wbs_dat_o[22]
port 391 nsew signal output
rlabel metal3 s 100 40992 400 41048 6 wbs_dat_o[23]
port 392 nsew signal output
rlabel metal2 s 26544 100 26600 400 6 wbs_dat_o[24]
port 393 nsew signal output
rlabel metal2 s 9408 100 9464 400 6 wbs_dat_o[25]
port 394 nsew signal output
rlabel metal2 s 64512 125592 64568 125892 6 wbs_dat_o[26]
port 395 nsew signal output
rlabel metal2 s 36624 125592 36680 125892 6 wbs_dat_o[27]
port 396 nsew signal output
rlabel metal2 s 67872 100 67928 400 6 wbs_dat_o[28]
port 397 nsew signal output
rlabel metal2 s 85344 125592 85400 125892 6 wbs_dat_o[29]
port 398 nsew signal output
rlabel metal3 s 123800 35952 124100 36008 6 wbs_dat_o[2]
port 399 nsew signal output
rlabel metal3 s 100 82320 400 82376 6 wbs_dat_o[30]
port 400 nsew signal output
rlabel metal3 s 123800 97776 124100 97832 6 wbs_dat_o[31]
port 401 nsew signal output
rlabel metal2 s 27888 100 27944 400 6 wbs_dat_o[3]
port 402 nsew signal output
rlabel metal2 s 48384 100 48440 400 6 wbs_dat_o[4]
port 403 nsew signal output
rlabel metal2 s 75264 100 75320 400 6 wbs_dat_o[5]
port 404 nsew signal output
rlabel metal3 s 123800 93072 124100 93128 6 wbs_dat_o[6]
port 405 nsew signal output
rlabel metal2 s 76272 100 76328 400 6 wbs_dat_o[7]
port 406 nsew signal output
rlabel metal2 s 81648 125592 81704 125892 6 wbs_dat_o[8]
port 407 nsew signal output
rlabel metal2 s 79296 125592 79352 125892 6 wbs_dat_o[9]
port 408 nsew signal output
rlabel metal3 s 100 115248 400 115304 6 wbs_sel_i[0]
port 409 nsew signal input
rlabel metal2 s 12432 125592 12488 125892 6 wbs_sel_i[1]
port 410 nsew signal input
rlabel metal2 s 91056 100 91112 400 6 wbs_sel_i[2]
port 411 nsew signal input
rlabel metal3 s 100 27888 400 27944 6 wbs_sel_i[3]
port 412 nsew signal input
rlabel metal3 s 100 103152 400 103208 6 wbs_stb_i
port 413 nsew signal input
rlabel metal3 s 123800 62496 124100 62552 6 wbs_we_i
port 414 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 124200 125992
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 41550244
string GDS_FILE /home/vijayan/CARAVEL_FLOW/GFmpw0/AES128_GFMPW0/openlane/aes_core/runs/22_12_03_09_58/results/signoff/aes_core.magic.gds
string GDS_START 335958
<< end >>

