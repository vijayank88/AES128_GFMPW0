VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aes_core
  CLASS BLOCK ;
  FOREIGN aes_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1154.760 BY 1172.680 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1168.680 679.280 1171.680 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 1168.680 148.400 1171.680 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 880.320 4.000 880.880 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1159.200 1153.760 1159.760 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.280 4.000 77.840 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 1168.680 850.640 1171.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 752.640 1153.760 753.200 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 540.960 4.000 541.520 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 423.360 1153.760 423.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1162.560 4.000 1163.120 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 1168.680 1132.880 1171.680 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 924.000 4.000 924.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 188.160 1153.760 188.720 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 598.080 4.000 598.640 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1168.680 249.200 1171.680 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1038.240 4.000 1038.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 1.000 995.120 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 245.280 1153.760 245.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 1.000 1129.520 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.760 4.000 54.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1142.400 1168.680 1142.960 1171.680 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 1168.680 588.560 1171.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.320 4.000 124.880 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 225.120 4.000 225.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 1168.680 554.960 1171.680 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1125.600 1153.760 1126.160 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1168.680 124.880 1171.680 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 876.960 1153.760 877.520 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 1168.680 985.040 1171.680 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 288.960 1153.760 289.520 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 406.560 4.000 407.120 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 493.920 1153.760 494.480 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 1168.680 91.280 1171.680 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 1168.680 941.360 1171.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 1.000 407.120 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 900.480 1153.760 901.040 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 1.000 235.760 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 107.520 1153.760 108.080 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 198.240 1153.760 198.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1.000 857.360 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1168.680 635.600 1171.680 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1128.960 4.000 1129.520 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 20.160 4.000 20.720 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1168.680 195.440 1171.680 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 1168.680 306.320 1171.680 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1168.680 158.480 1171.680 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 870.240 4.000 870.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 1.000 689.360 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1011.360 1153.760 1011.920 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 255.360 1153.760 255.920 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 890.400 4.000 890.960 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 1.000 1082.480 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1004.640 4.000 1005.200 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 1.000 958.160 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 1168.680 497.840 1171.680 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1168.680 622.160 1171.680 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1038.240 1.000 1038.800 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 413.280 1153.760 413.840 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 1168.680 837.200 1171.680 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 1168.680 974.960 1171.680 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 1.000 111.440 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1098.720 1168.680 1099.280 1171.680 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 1.000 460.880 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1168.680 171.920 1171.680 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 1168.680 47.600 1171.680 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 517.440 4.000 518.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 1.000 971.600 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 460.320 1153.760 460.880 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 1168.680 1018.640 1171.680 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 174.720 1153.760 175.280 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1065.120 1168.680 1065.680 1171.680 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1.000 484.400 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 1.000 722.960 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 131.040 1153.760 131.600 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 729.120 1153.760 729.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 789.600 4.000 790.160 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1058.400 1153.760 1058.960 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1168.680 521.360 1171.680 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1.000 134.960 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 779.520 4.000 780.080 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 1.000 746.480 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1.000 77.840 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 661.920 1153.760 662.480 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1.000 518.000 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 1.000 383.600 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 379.680 1153.760 380.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 1.000 981.680 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.760 4.000 474.320 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1085.280 1168.680 1085.840 1171.680 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1152.480 4.000 1153.040 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 608.160 4.000 608.720 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 766.080 1.000 766.640 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 1168.680 655.760 1171.680 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 732.480 4.000 733.040 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 231.840 1153.760 232.400 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 440.160 4.000 440.720 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 530.880 4.000 531.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 1.000 756.560 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 164.640 1153.760 165.200 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1149.120 1153.760 1149.680 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 40.320 1153.760 40.880 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1168.680 262.640 1171.680 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 1168.680 568.400 1171.680 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 483.840 4.000 484.400 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 675.360 4.000 675.920 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 1168.680 712.880 1171.680 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 1.000 833.840 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 1168.680 104.720 1171.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 349.440 4.000 350.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 1.000 1139.600 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1.000 427.280 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1.000 350.000 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 1168.680 477.680 1171.680 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 1168.680 1052.240 1171.680 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 1.000 541.520 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 708.960 4.000 709.520 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1168.680 904.400 1171.680 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1135.680 1153.760 1136.240 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 299.040 1153.760 299.600 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 756.000 4.000 756.560 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 221.760 1153.760 222.320 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 110.880 4.000 111.440 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 67.200 4.000 67.760 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 1168.680 927.920 1171.680 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 1168.680 726.320 1171.680 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 967.680 1153.760 968.240 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 1168.680 860.720 1171.680 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 564.480 4.000 565.040 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 994.560 4.000 995.120 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1068.480 1153.760 1069.040 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 638.400 1153.760 638.960 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1139.040 4.000 1139.600 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 480.480 1153.760 481.040 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1001.280 1153.760 1001.840 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 1.000 1095.920 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.800 4.000 269.360 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 1.000 813.680 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1168.680 420.560 1171.680 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 799.680 4.000 800.240 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 1168.680 487.760 1171.680 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 1168.680 780.080 1171.680 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 1.000 551.600 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1105.440 4.000 1106.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 497.280 4.000 497.840 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 823.200 4.000 823.760 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 843.360 1153.760 843.920 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 833.280 1153.760 833.840 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 100.800 4.000 101.360 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 87.360 4.000 87.920 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1.000 282.800 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1168.680 464.240 1171.680 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 1.000 531.440 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1061.760 4.000 1062.320 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 1168.680 353.360 1171.680 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 312.480 1153.760 313.040 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.840 4.000 316.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 325.920 4.000 326.480 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 30.240 1153.760 30.800 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 1.000 417.200 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 450.240 4.000 450.800 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 1.000 202.160 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 1168.680 803.600 1171.680 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 1168.680 884.240 1171.680 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 1.000 675.920 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 561.120 1153.760 561.680 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 574.560 4.000 575.120 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1168.680 0.560 1171.680 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 971.040 4.000 971.600 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1168.680 645.680 1171.680 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 168.000 4.000 168.560 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 722.400 4.000 722.960 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 1.000 823.760 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 846.720 4.000 847.280 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1168.680 329.840 1171.680 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 470.400 1153.760 470.960 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1092.000 1153.760 1092.560 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 628.320 1153.760 628.880 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 1168.680 578.480 1171.680 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1168.680 511.280 1171.680 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1.000 608.720 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 537.600 1153.760 538.160 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1168.680 544.880 1171.680 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 809.760 1153.760 810.320 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 1168.680 612.080 1171.680 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 178.080 4.000 178.640 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1.000 622.160 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1008.000 1168.680 1008.560 1171.680 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1.000 158.480 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 157.920 4.000 158.480 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 1.000 497.840 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 913.920 4.000 914.480 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 527.520 1153.760 528.080 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1168.680 34.160 1171.680 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1168.680 182.000 1171.680 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1168.680 24.080 1171.680 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1.000 565.040 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1.000 316.400 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 934.080 1153.760 934.640 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 446.880 1153.760 447.440 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 16.800 1153.760 17.360 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 154.560 1153.760 155.120 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 1168.680 817.040 1171.680 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1048.320 4.000 1048.880 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 346.080 1153.760 346.640 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 977.760 1153.760 978.320 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 1.000 67.760 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1.000 474.320 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 1168.680 702.800 1171.680 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1061.760 1.000 1062.320 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 833.280 4.000 833.840 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1.000 269.360 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1048.320 1.000 1048.880 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 1168.680 669.200 1171.680 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 1168.680 407.120 1171.680 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 426.720 4.000 427.280 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 73.920 1153.760 74.480 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 1.000 642.320 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1095.360 4.000 1095.920 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 1168.680 444.080 1171.680 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 265.440 1153.760 266.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 937.440 4.000 938.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 796.320 1153.760 796.880 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1034.880 1153.760 1035.440 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 695.520 1153.760 696.080 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 1168.680 951.440 1171.680 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 1.000 1005.200 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 87.360 1153.760 87.920 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 813.120 4.000 813.680 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 1168.680 1119.440 1171.680 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1081.920 4.000 1082.480 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 547.680 1153.760 548.240 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 436.800 1153.760 437.360 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 819.840 1153.760 820.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 651.840 1153.760 652.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 1168.680 454.160 1171.680 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 416.640 4.000 417.200 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.680 4.000 44.240 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 1.000 1015.280 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1.000 168.560 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.480 4.000 145.040 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 1168.680 81.200 1171.680 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 97.440 1153.760 98.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1168.680 229.040 1171.680 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1028.160 4.000 1028.720 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1168.680 205.520 1171.680 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.600 4.000 34.160 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 1.000 326.480 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 292.320 4.000 292.880 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 1.000 1028.720 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 1168.680 239.120 1171.680 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 1.000 212.240 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 604.800 1153.760 605.360 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1102.080 1153.760 1102.640 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 1168.680 1153.040 1171.680 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 991.200 1153.760 991.760 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 957.600 1153.760 958.160 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 944.160 1153.760 944.720 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 1.000 585.200 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1041.600 1168.680 1042.160 1171.680 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1.000 34.160 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 1.000 10.640 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 1168.680 14.000 1171.680 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1.000 598.640 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 507.360 4.000 507.920 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 641.760 4.000 642.320 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 372.960 4.000 373.520 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 1168.680 430.640 1171.680 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 745.920 4.000 746.480 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 1.000 225.680 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 1.000 507.920 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 584.640 4.000 585.200 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 1.000 924.560 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 1.000 440.720 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 856.800 4.000 857.360 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 571.200 1153.760 571.760 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 776.160 1153.760 776.720 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 1.000 890.960 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1168.680 373.520 1171.680 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 1.000 1153.040 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 742.560 1153.760 743.120 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 698.880 4.000 699.440 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 594.720 1153.760 595.280 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 1.000 880.880 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 1168.680 1028.720 1171.680 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 120.960 1153.760 121.520 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1168.680 692.720 1171.680 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 1.000 1072.400 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1168.680 282.800 1171.680 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1.000 145.040 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 10.080 4.000 10.640 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1118.880 4.000 1119.440 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 762.720 1153.760 763.280 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 1.000 292.880 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1105.440 1.000 1106.000 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 211.680 4.000 212.240 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 1168.680 995.120 1171.680 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 887.040 1153.760 887.600 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 1168.680 296.240 1171.680 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 1168.680 397.040 1171.680 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1156.700 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1156.700 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1156.700 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 211.680 1153.760 212.240 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 1168.680 215.600 1171.680 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 403.200 1153.760 403.760 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 1168.680 770.000 1171.680 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 1168.680 531.440 1171.680 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1168.680 71.120 1171.680 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 1.000 101.360 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 282.240 4.000 282.800 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 853.440 1153.760 854.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 786.240 1153.760 786.800 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 1.000 733.040 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 655.200 4.000 655.760 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 369.600 1153.760 370.160 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 1.000 1119.440 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 1168.680 746.480 1171.680 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 631.680 4.000 632.240 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 1.000 655.760 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 1.000 938.000 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 278.880 1153.760 279.440 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 1168.680 138.320 1171.680 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.600 4.000 202.160 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1.000 124.880 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1168.680 386.960 1171.680 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 685.440 1153.760 686.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1115.520 1153.760 1116.080 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.400 4.000 134.960 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 460.320 4.000 460.880 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 504.000 1153.760 504.560 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1.000 904.400 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 1168.680 894.320 1171.680 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 1.000 870.800 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1.000 373.520 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1.000 54.320 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 6.720 1153.760 7.280 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 322.560 1153.760 323.120 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1168.680 363.440 1171.680 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1024.800 1153.760 1025.360 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 903.840 4.000 904.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 981.120 4.000 981.680 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 947.520 4.000 948.080 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 1.000 44.240 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 618.240 1153.760 618.800 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.520 4.000 192.080 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1075.200 1168.680 1075.760 1171.680 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1168.680 57.680 1171.680 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1.000 178.640 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 708.960 1153.760 709.520 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1108.800 1168.680 1109.360 1171.680 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 688.800 4.000 689.360 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 920.640 1153.760 921.200 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 389.760 1153.760 390.320 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 1.000 800.240 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 1168.680 961.520 1171.680 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 1168.680 272.720 1171.680 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 1.000 360.080 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 719.040 1153.760 719.600 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 1.000 948.080 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 356.160 1153.760 356.720 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 621.600 4.000 622.160 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 50.400 1153.760 50.960 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1.000 192.080 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 1.000 575.120 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 514.080 1153.760 514.640 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 1168.680 917.840 1171.680 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1044.960 1153.760 1045.520 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 63.840 1153.760 64.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 235.200 4.000 235.760 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 672.000 1153.760 672.560 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 1.000 20.720 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 1081.920 1153.760 1082.480 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 1168.680 870.800 1171.680 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 141.120 1153.760 141.680 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 1168.680 827.120 1171.680 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1.000 790.160 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 359.520 4.000 360.080 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 1.000 780.080 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 1.000 914.480 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 551.040 4.000 551.600 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1014.720 4.000 1015.280 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 1168.680 319.760 1171.680 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 383.040 4.000 383.600 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 1.000 87.920 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 1168.680 602.000 1171.680 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 1168.680 339.920 1171.680 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 1.000 632.240 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 1168.680 793.520 1171.680 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 336.000 1153.760 336.560 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 766.080 4.000 766.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 910.560 1153.760 911.120 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1.000 259.280 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 1.000 450.800 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 1.000 699.440 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 866.880 1153.760 867.440 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 1.000 709.520 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1168.680 759.920 1171.680 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 1168.680 736.400 1171.680 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1071.840 4.000 1072.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1168.680 114.800 1171.680 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 1.000 847.280 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.720 4.000 259.280 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 957.600 4.000 958.160 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1150.760 584.640 1153.760 585.200 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 1148.000 1157.370 ;
      LAYER Metal2 ;
        RECT 0.860 1168.380 13.140 1169.140 ;
        RECT 14.300 1168.380 23.220 1169.140 ;
        RECT 24.380 1168.380 33.300 1169.140 ;
        RECT 34.460 1168.380 46.740 1169.140 ;
        RECT 47.900 1168.380 56.820 1169.140 ;
        RECT 57.980 1168.380 70.260 1169.140 ;
        RECT 71.420 1168.380 80.340 1169.140 ;
        RECT 81.500 1168.380 90.420 1169.140 ;
        RECT 91.580 1168.380 103.860 1169.140 ;
        RECT 105.020 1168.380 113.940 1169.140 ;
        RECT 115.100 1168.380 124.020 1169.140 ;
        RECT 125.180 1168.380 137.460 1169.140 ;
        RECT 138.620 1168.380 147.540 1169.140 ;
        RECT 148.700 1168.380 157.620 1169.140 ;
        RECT 158.780 1168.380 171.060 1169.140 ;
        RECT 172.220 1168.380 181.140 1169.140 ;
        RECT 182.300 1168.380 194.580 1169.140 ;
        RECT 195.740 1168.380 204.660 1169.140 ;
        RECT 205.820 1168.380 214.740 1169.140 ;
        RECT 215.900 1168.380 228.180 1169.140 ;
        RECT 229.340 1168.380 238.260 1169.140 ;
        RECT 239.420 1168.380 248.340 1169.140 ;
        RECT 249.500 1168.380 261.780 1169.140 ;
        RECT 262.940 1168.380 271.860 1169.140 ;
        RECT 273.020 1168.380 281.940 1169.140 ;
        RECT 283.100 1168.380 295.380 1169.140 ;
        RECT 296.540 1168.380 305.460 1169.140 ;
        RECT 306.620 1168.380 318.900 1169.140 ;
        RECT 320.060 1168.380 328.980 1169.140 ;
        RECT 330.140 1168.380 339.060 1169.140 ;
        RECT 340.220 1168.380 352.500 1169.140 ;
        RECT 353.660 1168.380 362.580 1169.140 ;
        RECT 363.740 1168.380 372.660 1169.140 ;
        RECT 373.820 1168.380 386.100 1169.140 ;
        RECT 387.260 1168.380 396.180 1169.140 ;
        RECT 397.340 1168.380 406.260 1169.140 ;
        RECT 407.420 1168.380 419.700 1169.140 ;
        RECT 420.860 1168.380 429.780 1169.140 ;
        RECT 430.940 1168.380 443.220 1169.140 ;
        RECT 444.380 1168.380 453.300 1169.140 ;
        RECT 454.460 1168.380 463.380 1169.140 ;
        RECT 464.540 1168.380 476.820 1169.140 ;
        RECT 477.980 1168.380 486.900 1169.140 ;
        RECT 488.060 1168.380 496.980 1169.140 ;
        RECT 498.140 1168.380 510.420 1169.140 ;
        RECT 511.580 1168.380 520.500 1169.140 ;
        RECT 521.660 1168.380 530.580 1169.140 ;
        RECT 531.740 1168.380 544.020 1169.140 ;
        RECT 545.180 1168.380 554.100 1169.140 ;
        RECT 555.260 1168.380 567.540 1169.140 ;
        RECT 568.700 1168.380 577.620 1169.140 ;
        RECT 578.780 1168.380 587.700 1169.140 ;
        RECT 588.860 1168.380 601.140 1169.140 ;
        RECT 602.300 1168.380 611.220 1169.140 ;
        RECT 612.380 1168.380 621.300 1169.140 ;
        RECT 622.460 1168.380 634.740 1169.140 ;
        RECT 635.900 1168.380 644.820 1169.140 ;
        RECT 645.980 1168.380 654.900 1169.140 ;
        RECT 656.060 1168.380 668.340 1169.140 ;
        RECT 669.500 1168.380 678.420 1169.140 ;
        RECT 679.580 1168.380 691.860 1169.140 ;
        RECT 693.020 1168.380 701.940 1169.140 ;
        RECT 703.100 1168.380 712.020 1169.140 ;
        RECT 713.180 1168.380 725.460 1169.140 ;
        RECT 726.620 1168.380 735.540 1169.140 ;
        RECT 736.700 1168.380 745.620 1169.140 ;
        RECT 746.780 1168.380 759.060 1169.140 ;
        RECT 760.220 1168.380 769.140 1169.140 ;
        RECT 770.300 1168.380 779.220 1169.140 ;
        RECT 780.380 1168.380 792.660 1169.140 ;
        RECT 793.820 1168.380 802.740 1169.140 ;
        RECT 803.900 1168.380 816.180 1169.140 ;
        RECT 817.340 1168.380 826.260 1169.140 ;
        RECT 827.420 1168.380 836.340 1169.140 ;
        RECT 837.500 1168.380 849.780 1169.140 ;
        RECT 850.940 1168.380 859.860 1169.140 ;
        RECT 861.020 1168.380 869.940 1169.140 ;
        RECT 871.100 1168.380 883.380 1169.140 ;
        RECT 884.540 1168.380 893.460 1169.140 ;
        RECT 894.620 1168.380 903.540 1169.140 ;
        RECT 904.700 1168.380 916.980 1169.140 ;
        RECT 918.140 1168.380 927.060 1169.140 ;
        RECT 928.220 1168.380 940.500 1169.140 ;
        RECT 941.660 1168.380 950.580 1169.140 ;
        RECT 951.740 1168.380 960.660 1169.140 ;
        RECT 961.820 1168.380 974.100 1169.140 ;
        RECT 975.260 1168.380 984.180 1169.140 ;
        RECT 985.340 1168.380 994.260 1169.140 ;
        RECT 995.420 1168.380 1007.700 1169.140 ;
        RECT 1008.860 1168.380 1017.780 1169.140 ;
        RECT 1018.940 1168.380 1027.860 1169.140 ;
        RECT 1029.020 1168.380 1041.300 1169.140 ;
        RECT 1042.460 1168.380 1051.380 1169.140 ;
        RECT 1052.540 1168.380 1064.820 1169.140 ;
        RECT 1065.980 1168.380 1074.900 1169.140 ;
        RECT 1076.060 1168.380 1084.980 1169.140 ;
        RECT 1086.140 1168.380 1098.420 1169.140 ;
        RECT 1099.580 1168.380 1108.500 1169.140 ;
        RECT 1109.660 1168.380 1118.580 1169.140 ;
        RECT 1119.740 1168.380 1132.020 1169.140 ;
        RECT 1133.180 1168.380 1142.100 1169.140 ;
        RECT 1143.260 1168.380 1146.740 1169.140 ;
        RECT 0.140 4.300 1146.740 1168.380 ;
        RECT 0.860 4.000 9.780 4.300 ;
        RECT 10.940 4.000 19.860 4.300 ;
        RECT 21.020 4.000 33.300 4.300 ;
        RECT 34.460 4.000 43.380 4.300 ;
        RECT 44.540 4.000 53.460 4.300 ;
        RECT 54.620 4.000 66.900 4.300 ;
        RECT 68.060 4.000 76.980 4.300 ;
        RECT 78.140 4.000 87.060 4.300 ;
        RECT 88.220 4.000 100.500 4.300 ;
        RECT 101.660 4.000 110.580 4.300 ;
        RECT 111.740 4.000 124.020 4.300 ;
        RECT 125.180 4.000 134.100 4.300 ;
        RECT 135.260 4.000 144.180 4.300 ;
        RECT 145.340 4.000 157.620 4.300 ;
        RECT 158.780 4.000 167.700 4.300 ;
        RECT 168.860 4.000 177.780 4.300 ;
        RECT 178.940 4.000 191.220 4.300 ;
        RECT 192.380 4.000 201.300 4.300 ;
        RECT 202.460 4.000 211.380 4.300 ;
        RECT 212.540 4.000 224.820 4.300 ;
        RECT 225.980 4.000 234.900 4.300 ;
        RECT 236.060 4.000 248.340 4.300 ;
        RECT 249.500 4.000 258.420 4.300 ;
        RECT 259.580 4.000 268.500 4.300 ;
        RECT 269.660 4.000 281.940 4.300 ;
        RECT 283.100 4.000 292.020 4.300 ;
        RECT 293.180 4.000 302.100 4.300 ;
        RECT 303.260 4.000 315.540 4.300 ;
        RECT 316.700 4.000 325.620 4.300 ;
        RECT 326.780 4.000 335.700 4.300 ;
        RECT 336.860 4.000 349.140 4.300 ;
        RECT 350.300 4.000 359.220 4.300 ;
        RECT 360.380 4.000 372.660 4.300 ;
        RECT 373.820 4.000 382.740 4.300 ;
        RECT 383.900 4.000 392.820 4.300 ;
        RECT 393.980 4.000 406.260 4.300 ;
        RECT 407.420 4.000 416.340 4.300 ;
        RECT 417.500 4.000 426.420 4.300 ;
        RECT 427.580 4.000 439.860 4.300 ;
        RECT 441.020 4.000 449.940 4.300 ;
        RECT 451.100 4.000 460.020 4.300 ;
        RECT 461.180 4.000 473.460 4.300 ;
        RECT 474.620 4.000 483.540 4.300 ;
        RECT 484.700 4.000 496.980 4.300 ;
        RECT 498.140 4.000 507.060 4.300 ;
        RECT 508.220 4.000 517.140 4.300 ;
        RECT 518.300 4.000 530.580 4.300 ;
        RECT 531.740 4.000 540.660 4.300 ;
        RECT 541.820 4.000 550.740 4.300 ;
        RECT 551.900 4.000 564.180 4.300 ;
        RECT 565.340 4.000 574.260 4.300 ;
        RECT 575.420 4.000 584.340 4.300 ;
        RECT 585.500 4.000 597.780 4.300 ;
        RECT 598.940 4.000 607.860 4.300 ;
        RECT 609.020 4.000 621.300 4.300 ;
        RECT 622.460 4.000 631.380 4.300 ;
        RECT 632.540 4.000 641.460 4.300 ;
        RECT 642.620 4.000 654.900 4.300 ;
        RECT 656.060 4.000 664.980 4.300 ;
        RECT 666.140 4.000 675.060 4.300 ;
        RECT 676.220 4.000 688.500 4.300 ;
        RECT 689.660 4.000 698.580 4.300 ;
        RECT 699.740 4.000 708.660 4.300 ;
        RECT 709.820 4.000 722.100 4.300 ;
        RECT 723.260 4.000 732.180 4.300 ;
        RECT 733.340 4.000 745.620 4.300 ;
        RECT 746.780 4.000 755.700 4.300 ;
        RECT 756.860 4.000 765.780 4.300 ;
        RECT 766.940 4.000 779.220 4.300 ;
        RECT 780.380 4.000 789.300 4.300 ;
        RECT 790.460 4.000 799.380 4.300 ;
        RECT 800.540 4.000 812.820 4.300 ;
        RECT 813.980 4.000 822.900 4.300 ;
        RECT 824.060 4.000 832.980 4.300 ;
        RECT 834.140 4.000 846.420 4.300 ;
        RECT 847.580 4.000 856.500 4.300 ;
        RECT 857.660 4.000 869.940 4.300 ;
        RECT 871.100 4.000 880.020 4.300 ;
        RECT 881.180 4.000 890.100 4.300 ;
        RECT 891.260 4.000 903.540 4.300 ;
        RECT 904.700 4.000 913.620 4.300 ;
        RECT 914.780 4.000 923.700 4.300 ;
        RECT 924.860 4.000 937.140 4.300 ;
        RECT 938.300 4.000 947.220 4.300 ;
        RECT 948.380 4.000 957.300 4.300 ;
        RECT 958.460 4.000 970.740 4.300 ;
        RECT 971.900 4.000 980.820 4.300 ;
        RECT 981.980 4.000 994.260 4.300 ;
        RECT 995.420 4.000 1004.340 4.300 ;
        RECT 1005.500 4.000 1014.420 4.300 ;
        RECT 1015.580 4.000 1027.860 4.300 ;
        RECT 1029.020 4.000 1037.940 4.300 ;
        RECT 1039.100 4.000 1048.020 4.300 ;
        RECT 1049.180 4.000 1061.460 4.300 ;
        RECT 1062.620 4.000 1071.540 4.300 ;
        RECT 1072.700 4.000 1081.620 4.300 ;
        RECT 1082.780 4.000 1095.060 4.300 ;
        RECT 1096.220 4.000 1105.140 4.300 ;
        RECT 1106.300 4.000 1118.580 4.300 ;
        RECT 1119.740 4.000 1128.660 4.300 ;
        RECT 1129.820 4.000 1138.740 4.300 ;
        RECT 1139.900 4.000 1146.740 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 1153.340 1150.760 1157.380 ;
        RECT 0.090 1152.180 0.700 1153.340 ;
        RECT 4.300 1152.180 1150.760 1153.340 ;
        RECT 0.090 1149.980 1150.760 1152.180 ;
        RECT 0.090 1148.820 1150.460 1149.980 ;
        RECT 0.090 1139.900 1150.760 1148.820 ;
        RECT 0.090 1138.740 0.700 1139.900 ;
        RECT 4.300 1138.740 1150.760 1139.900 ;
        RECT 0.090 1136.540 1150.760 1138.740 ;
        RECT 0.090 1135.380 1150.460 1136.540 ;
        RECT 0.090 1129.820 1150.760 1135.380 ;
        RECT 0.090 1128.660 0.700 1129.820 ;
        RECT 4.300 1128.660 1150.760 1129.820 ;
        RECT 0.090 1126.460 1150.760 1128.660 ;
        RECT 0.090 1125.300 1150.460 1126.460 ;
        RECT 0.090 1119.740 1150.760 1125.300 ;
        RECT 0.090 1118.580 0.700 1119.740 ;
        RECT 4.300 1118.580 1150.760 1119.740 ;
        RECT 0.090 1116.380 1150.760 1118.580 ;
        RECT 0.090 1115.220 1150.460 1116.380 ;
        RECT 0.090 1106.300 1150.760 1115.220 ;
        RECT 0.090 1105.140 0.700 1106.300 ;
        RECT 4.300 1105.140 1150.760 1106.300 ;
        RECT 0.090 1102.940 1150.760 1105.140 ;
        RECT 0.090 1101.780 1150.460 1102.940 ;
        RECT 0.090 1096.220 1150.760 1101.780 ;
        RECT 0.090 1095.060 0.700 1096.220 ;
        RECT 4.300 1095.060 1150.760 1096.220 ;
        RECT 0.090 1092.860 1150.760 1095.060 ;
        RECT 0.090 1091.700 1150.460 1092.860 ;
        RECT 0.090 1082.780 1150.760 1091.700 ;
        RECT 0.090 1081.620 0.700 1082.780 ;
        RECT 4.300 1081.620 1150.460 1082.780 ;
        RECT 0.090 1072.700 1150.760 1081.620 ;
        RECT 0.090 1071.540 0.700 1072.700 ;
        RECT 4.300 1071.540 1150.760 1072.700 ;
        RECT 0.090 1069.340 1150.760 1071.540 ;
        RECT 0.090 1068.180 1150.460 1069.340 ;
        RECT 0.090 1062.620 1150.760 1068.180 ;
        RECT 0.090 1061.460 0.700 1062.620 ;
        RECT 4.300 1061.460 1150.760 1062.620 ;
        RECT 0.090 1059.260 1150.760 1061.460 ;
        RECT 0.090 1058.100 1150.460 1059.260 ;
        RECT 0.090 1049.180 1150.760 1058.100 ;
        RECT 0.090 1048.020 0.700 1049.180 ;
        RECT 4.300 1048.020 1150.760 1049.180 ;
        RECT 0.090 1045.820 1150.760 1048.020 ;
        RECT 0.090 1044.660 1150.460 1045.820 ;
        RECT 0.090 1039.100 1150.760 1044.660 ;
        RECT 0.090 1037.940 0.700 1039.100 ;
        RECT 4.300 1037.940 1150.760 1039.100 ;
        RECT 0.090 1035.740 1150.760 1037.940 ;
        RECT 0.090 1034.580 1150.460 1035.740 ;
        RECT 0.090 1029.020 1150.760 1034.580 ;
        RECT 0.090 1027.860 0.700 1029.020 ;
        RECT 4.300 1027.860 1150.760 1029.020 ;
        RECT 0.090 1025.660 1150.760 1027.860 ;
        RECT 0.090 1024.500 1150.460 1025.660 ;
        RECT 0.090 1015.580 1150.760 1024.500 ;
        RECT 0.090 1014.420 0.700 1015.580 ;
        RECT 4.300 1014.420 1150.760 1015.580 ;
        RECT 0.090 1012.220 1150.760 1014.420 ;
        RECT 0.090 1011.060 1150.460 1012.220 ;
        RECT 0.090 1005.500 1150.760 1011.060 ;
        RECT 0.090 1004.340 0.700 1005.500 ;
        RECT 4.300 1004.340 1150.760 1005.500 ;
        RECT 0.090 1002.140 1150.760 1004.340 ;
        RECT 0.090 1000.980 1150.460 1002.140 ;
        RECT 0.090 995.420 1150.760 1000.980 ;
        RECT 0.090 994.260 0.700 995.420 ;
        RECT 4.300 994.260 1150.760 995.420 ;
        RECT 0.090 992.060 1150.760 994.260 ;
        RECT 0.090 990.900 1150.460 992.060 ;
        RECT 0.090 981.980 1150.760 990.900 ;
        RECT 0.090 980.820 0.700 981.980 ;
        RECT 4.300 980.820 1150.760 981.980 ;
        RECT 0.090 978.620 1150.760 980.820 ;
        RECT 0.090 977.460 1150.460 978.620 ;
        RECT 0.090 971.900 1150.760 977.460 ;
        RECT 0.090 970.740 0.700 971.900 ;
        RECT 4.300 970.740 1150.760 971.900 ;
        RECT 0.090 968.540 1150.760 970.740 ;
        RECT 0.090 967.380 1150.460 968.540 ;
        RECT 0.090 958.460 1150.760 967.380 ;
        RECT 0.090 957.300 0.700 958.460 ;
        RECT 4.300 957.300 1150.460 958.460 ;
        RECT 0.090 948.380 1150.760 957.300 ;
        RECT 0.090 947.220 0.700 948.380 ;
        RECT 4.300 947.220 1150.760 948.380 ;
        RECT 0.090 945.020 1150.760 947.220 ;
        RECT 0.090 943.860 1150.460 945.020 ;
        RECT 0.090 938.300 1150.760 943.860 ;
        RECT 0.090 937.140 0.700 938.300 ;
        RECT 4.300 937.140 1150.760 938.300 ;
        RECT 0.090 934.940 1150.760 937.140 ;
        RECT 0.090 933.780 1150.460 934.940 ;
        RECT 0.090 924.860 1150.760 933.780 ;
        RECT 0.090 923.700 0.700 924.860 ;
        RECT 4.300 923.700 1150.760 924.860 ;
        RECT 0.090 921.500 1150.760 923.700 ;
        RECT 0.090 920.340 1150.460 921.500 ;
        RECT 0.090 914.780 1150.760 920.340 ;
        RECT 0.090 913.620 0.700 914.780 ;
        RECT 4.300 913.620 1150.760 914.780 ;
        RECT 0.090 911.420 1150.760 913.620 ;
        RECT 0.090 910.260 1150.460 911.420 ;
        RECT 0.090 904.700 1150.760 910.260 ;
        RECT 0.090 903.540 0.700 904.700 ;
        RECT 4.300 903.540 1150.760 904.700 ;
        RECT 0.090 901.340 1150.760 903.540 ;
        RECT 0.090 900.180 1150.460 901.340 ;
        RECT 0.090 891.260 1150.760 900.180 ;
        RECT 0.090 890.100 0.700 891.260 ;
        RECT 4.300 890.100 1150.760 891.260 ;
        RECT 0.090 887.900 1150.760 890.100 ;
        RECT 0.090 886.740 1150.460 887.900 ;
        RECT 0.090 881.180 1150.760 886.740 ;
        RECT 0.090 880.020 0.700 881.180 ;
        RECT 4.300 880.020 1150.760 881.180 ;
        RECT 0.090 877.820 1150.760 880.020 ;
        RECT 0.090 876.660 1150.460 877.820 ;
        RECT 0.090 871.100 1150.760 876.660 ;
        RECT 0.090 869.940 0.700 871.100 ;
        RECT 4.300 869.940 1150.760 871.100 ;
        RECT 0.090 867.740 1150.760 869.940 ;
        RECT 0.090 866.580 1150.460 867.740 ;
        RECT 0.090 857.660 1150.760 866.580 ;
        RECT 0.090 856.500 0.700 857.660 ;
        RECT 4.300 856.500 1150.760 857.660 ;
        RECT 0.090 854.300 1150.760 856.500 ;
        RECT 0.090 853.140 1150.460 854.300 ;
        RECT 0.090 847.580 1150.760 853.140 ;
        RECT 0.090 846.420 0.700 847.580 ;
        RECT 4.300 846.420 1150.760 847.580 ;
        RECT 0.090 844.220 1150.760 846.420 ;
        RECT 0.090 843.060 1150.460 844.220 ;
        RECT 0.090 834.140 1150.760 843.060 ;
        RECT 0.090 832.980 0.700 834.140 ;
        RECT 4.300 832.980 1150.460 834.140 ;
        RECT 0.090 824.060 1150.760 832.980 ;
        RECT 0.090 822.900 0.700 824.060 ;
        RECT 4.300 822.900 1150.760 824.060 ;
        RECT 0.090 820.700 1150.760 822.900 ;
        RECT 0.090 819.540 1150.460 820.700 ;
        RECT 0.090 813.980 1150.760 819.540 ;
        RECT 0.090 812.820 0.700 813.980 ;
        RECT 4.300 812.820 1150.760 813.980 ;
        RECT 0.090 810.620 1150.760 812.820 ;
        RECT 0.090 809.460 1150.460 810.620 ;
        RECT 0.090 800.540 1150.760 809.460 ;
        RECT 0.090 799.380 0.700 800.540 ;
        RECT 4.300 799.380 1150.760 800.540 ;
        RECT 0.090 797.180 1150.760 799.380 ;
        RECT 0.090 796.020 1150.460 797.180 ;
        RECT 0.090 790.460 1150.760 796.020 ;
        RECT 0.090 789.300 0.700 790.460 ;
        RECT 4.300 789.300 1150.760 790.460 ;
        RECT 0.090 787.100 1150.760 789.300 ;
        RECT 0.090 785.940 1150.460 787.100 ;
        RECT 0.090 780.380 1150.760 785.940 ;
        RECT 0.090 779.220 0.700 780.380 ;
        RECT 4.300 779.220 1150.760 780.380 ;
        RECT 0.090 777.020 1150.760 779.220 ;
        RECT 0.090 775.860 1150.460 777.020 ;
        RECT 0.090 766.940 1150.760 775.860 ;
        RECT 0.090 765.780 0.700 766.940 ;
        RECT 4.300 765.780 1150.760 766.940 ;
        RECT 0.090 763.580 1150.760 765.780 ;
        RECT 0.090 762.420 1150.460 763.580 ;
        RECT 0.090 756.860 1150.760 762.420 ;
        RECT 0.090 755.700 0.700 756.860 ;
        RECT 4.300 755.700 1150.760 756.860 ;
        RECT 0.090 753.500 1150.760 755.700 ;
        RECT 0.090 752.340 1150.460 753.500 ;
        RECT 0.090 746.780 1150.760 752.340 ;
        RECT 0.090 745.620 0.700 746.780 ;
        RECT 4.300 745.620 1150.760 746.780 ;
        RECT 0.090 743.420 1150.760 745.620 ;
        RECT 0.090 742.260 1150.460 743.420 ;
        RECT 0.090 733.340 1150.760 742.260 ;
        RECT 0.090 732.180 0.700 733.340 ;
        RECT 4.300 732.180 1150.760 733.340 ;
        RECT 0.090 729.980 1150.760 732.180 ;
        RECT 0.090 728.820 1150.460 729.980 ;
        RECT 0.090 723.260 1150.760 728.820 ;
        RECT 0.090 722.100 0.700 723.260 ;
        RECT 4.300 722.100 1150.760 723.260 ;
        RECT 0.090 719.900 1150.760 722.100 ;
        RECT 0.090 718.740 1150.460 719.900 ;
        RECT 0.090 709.820 1150.760 718.740 ;
        RECT 0.090 708.660 0.700 709.820 ;
        RECT 4.300 708.660 1150.460 709.820 ;
        RECT 0.090 699.740 1150.760 708.660 ;
        RECT 0.090 698.580 0.700 699.740 ;
        RECT 4.300 698.580 1150.760 699.740 ;
        RECT 0.090 696.380 1150.760 698.580 ;
        RECT 0.090 695.220 1150.460 696.380 ;
        RECT 0.090 689.660 1150.760 695.220 ;
        RECT 0.090 688.500 0.700 689.660 ;
        RECT 4.300 688.500 1150.760 689.660 ;
        RECT 0.090 686.300 1150.760 688.500 ;
        RECT 0.090 685.140 1150.460 686.300 ;
        RECT 0.090 676.220 1150.760 685.140 ;
        RECT 0.090 675.060 0.700 676.220 ;
        RECT 4.300 675.060 1150.760 676.220 ;
        RECT 0.090 672.860 1150.760 675.060 ;
        RECT 0.090 671.700 1150.460 672.860 ;
        RECT 0.090 666.140 1150.760 671.700 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 1150.760 666.140 ;
        RECT 0.090 662.780 1150.760 664.980 ;
        RECT 0.090 661.620 1150.460 662.780 ;
        RECT 0.090 656.060 1150.760 661.620 ;
        RECT 0.090 654.900 0.700 656.060 ;
        RECT 4.300 654.900 1150.760 656.060 ;
        RECT 0.090 652.700 1150.760 654.900 ;
        RECT 0.090 651.540 1150.460 652.700 ;
        RECT 0.090 642.620 1150.760 651.540 ;
        RECT 0.090 641.460 0.700 642.620 ;
        RECT 4.300 641.460 1150.760 642.620 ;
        RECT 0.090 639.260 1150.760 641.460 ;
        RECT 0.090 638.100 1150.460 639.260 ;
        RECT 0.090 632.540 1150.760 638.100 ;
        RECT 0.090 631.380 0.700 632.540 ;
        RECT 4.300 631.380 1150.760 632.540 ;
        RECT 0.090 629.180 1150.760 631.380 ;
        RECT 0.090 628.020 1150.460 629.180 ;
        RECT 0.090 622.460 1150.760 628.020 ;
        RECT 0.090 621.300 0.700 622.460 ;
        RECT 4.300 621.300 1150.760 622.460 ;
        RECT 0.090 619.100 1150.760 621.300 ;
        RECT 0.090 617.940 1150.460 619.100 ;
        RECT 0.090 609.020 1150.760 617.940 ;
        RECT 0.090 607.860 0.700 609.020 ;
        RECT 4.300 607.860 1150.760 609.020 ;
        RECT 0.090 605.660 1150.760 607.860 ;
        RECT 0.090 604.500 1150.460 605.660 ;
        RECT 0.090 598.940 1150.760 604.500 ;
        RECT 0.090 597.780 0.700 598.940 ;
        RECT 4.300 597.780 1150.760 598.940 ;
        RECT 0.090 595.580 1150.760 597.780 ;
        RECT 0.090 594.420 1150.460 595.580 ;
        RECT 0.090 585.500 1150.760 594.420 ;
        RECT 0.090 584.340 0.700 585.500 ;
        RECT 4.300 584.340 1150.460 585.500 ;
        RECT 0.090 575.420 1150.760 584.340 ;
        RECT 0.090 574.260 0.700 575.420 ;
        RECT 4.300 574.260 1150.760 575.420 ;
        RECT 0.090 572.060 1150.760 574.260 ;
        RECT 0.090 570.900 1150.460 572.060 ;
        RECT 0.090 565.340 1150.760 570.900 ;
        RECT 0.090 564.180 0.700 565.340 ;
        RECT 4.300 564.180 1150.760 565.340 ;
        RECT 0.090 561.980 1150.760 564.180 ;
        RECT 0.090 560.820 1150.460 561.980 ;
        RECT 0.090 551.900 1150.760 560.820 ;
        RECT 0.090 550.740 0.700 551.900 ;
        RECT 4.300 550.740 1150.760 551.900 ;
        RECT 0.090 548.540 1150.760 550.740 ;
        RECT 0.090 547.380 1150.460 548.540 ;
        RECT 0.090 541.820 1150.760 547.380 ;
        RECT 0.090 540.660 0.700 541.820 ;
        RECT 4.300 540.660 1150.760 541.820 ;
        RECT 0.090 538.460 1150.760 540.660 ;
        RECT 0.090 537.300 1150.460 538.460 ;
        RECT 0.090 531.740 1150.760 537.300 ;
        RECT 0.090 530.580 0.700 531.740 ;
        RECT 4.300 530.580 1150.760 531.740 ;
        RECT 0.090 528.380 1150.760 530.580 ;
        RECT 0.090 527.220 1150.460 528.380 ;
        RECT 0.090 518.300 1150.760 527.220 ;
        RECT 0.090 517.140 0.700 518.300 ;
        RECT 4.300 517.140 1150.760 518.300 ;
        RECT 0.090 514.940 1150.760 517.140 ;
        RECT 0.090 513.780 1150.460 514.940 ;
        RECT 0.090 508.220 1150.760 513.780 ;
        RECT 0.090 507.060 0.700 508.220 ;
        RECT 4.300 507.060 1150.760 508.220 ;
        RECT 0.090 504.860 1150.760 507.060 ;
        RECT 0.090 503.700 1150.460 504.860 ;
        RECT 0.090 498.140 1150.760 503.700 ;
        RECT 0.090 496.980 0.700 498.140 ;
        RECT 4.300 496.980 1150.760 498.140 ;
        RECT 0.090 494.780 1150.760 496.980 ;
        RECT 0.090 493.620 1150.460 494.780 ;
        RECT 0.090 484.700 1150.760 493.620 ;
        RECT 0.090 483.540 0.700 484.700 ;
        RECT 4.300 483.540 1150.760 484.700 ;
        RECT 0.090 481.340 1150.760 483.540 ;
        RECT 0.090 480.180 1150.460 481.340 ;
        RECT 0.090 474.620 1150.760 480.180 ;
        RECT 0.090 473.460 0.700 474.620 ;
        RECT 4.300 473.460 1150.760 474.620 ;
        RECT 0.090 471.260 1150.760 473.460 ;
        RECT 0.090 470.100 1150.460 471.260 ;
        RECT 0.090 461.180 1150.760 470.100 ;
        RECT 0.090 460.020 0.700 461.180 ;
        RECT 4.300 460.020 1150.460 461.180 ;
        RECT 0.090 451.100 1150.760 460.020 ;
        RECT 0.090 449.940 0.700 451.100 ;
        RECT 4.300 449.940 1150.760 451.100 ;
        RECT 0.090 447.740 1150.760 449.940 ;
        RECT 0.090 446.580 1150.460 447.740 ;
        RECT 0.090 441.020 1150.760 446.580 ;
        RECT 0.090 439.860 0.700 441.020 ;
        RECT 4.300 439.860 1150.760 441.020 ;
        RECT 0.090 437.660 1150.760 439.860 ;
        RECT 0.090 436.500 1150.460 437.660 ;
        RECT 0.090 427.580 1150.760 436.500 ;
        RECT 0.090 426.420 0.700 427.580 ;
        RECT 4.300 426.420 1150.760 427.580 ;
        RECT 0.090 424.220 1150.760 426.420 ;
        RECT 0.090 423.060 1150.460 424.220 ;
        RECT 0.090 417.500 1150.760 423.060 ;
        RECT 0.090 416.340 0.700 417.500 ;
        RECT 4.300 416.340 1150.760 417.500 ;
        RECT 0.090 414.140 1150.760 416.340 ;
        RECT 0.090 412.980 1150.460 414.140 ;
        RECT 0.090 407.420 1150.760 412.980 ;
        RECT 0.090 406.260 0.700 407.420 ;
        RECT 4.300 406.260 1150.760 407.420 ;
        RECT 0.090 404.060 1150.760 406.260 ;
        RECT 0.090 402.900 1150.460 404.060 ;
        RECT 0.090 393.980 1150.760 402.900 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 1150.760 393.980 ;
        RECT 0.090 390.620 1150.760 392.820 ;
        RECT 0.090 389.460 1150.460 390.620 ;
        RECT 0.090 383.900 1150.760 389.460 ;
        RECT 0.090 382.740 0.700 383.900 ;
        RECT 4.300 382.740 1150.760 383.900 ;
        RECT 0.090 380.540 1150.760 382.740 ;
        RECT 0.090 379.380 1150.460 380.540 ;
        RECT 0.090 373.820 1150.760 379.380 ;
        RECT 0.090 372.660 0.700 373.820 ;
        RECT 4.300 372.660 1150.760 373.820 ;
        RECT 0.090 370.460 1150.760 372.660 ;
        RECT 0.090 369.300 1150.460 370.460 ;
        RECT 0.090 360.380 1150.760 369.300 ;
        RECT 0.090 359.220 0.700 360.380 ;
        RECT 4.300 359.220 1150.760 360.380 ;
        RECT 0.090 357.020 1150.760 359.220 ;
        RECT 0.090 355.860 1150.460 357.020 ;
        RECT 0.090 350.300 1150.760 355.860 ;
        RECT 0.090 349.140 0.700 350.300 ;
        RECT 4.300 349.140 1150.760 350.300 ;
        RECT 0.090 346.940 1150.760 349.140 ;
        RECT 0.090 345.780 1150.460 346.940 ;
        RECT 0.090 336.860 1150.760 345.780 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 1150.460 336.860 ;
        RECT 0.090 326.780 1150.760 335.700 ;
        RECT 0.090 325.620 0.700 326.780 ;
        RECT 4.300 325.620 1150.760 326.780 ;
        RECT 0.090 323.420 1150.760 325.620 ;
        RECT 0.090 322.260 1150.460 323.420 ;
        RECT 0.090 316.700 1150.760 322.260 ;
        RECT 0.090 315.540 0.700 316.700 ;
        RECT 4.300 315.540 1150.760 316.700 ;
        RECT 0.090 313.340 1150.760 315.540 ;
        RECT 0.090 312.180 1150.460 313.340 ;
        RECT 0.090 303.260 1150.760 312.180 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 1150.760 303.260 ;
        RECT 0.090 299.900 1150.760 302.100 ;
        RECT 0.090 298.740 1150.460 299.900 ;
        RECT 0.090 293.180 1150.760 298.740 ;
        RECT 0.090 292.020 0.700 293.180 ;
        RECT 4.300 292.020 1150.760 293.180 ;
        RECT 0.090 289.820 1150.760 292.020 ;
        RECT 0.090 288.660 1150.460 289.820 ;
        RECT 0.090 283.100 1150.760 288.660 ;
        RECT 0.090 281.940 0.700 283.100 ;
        RECT 4.300 281.940 1150.760 283.100 ;
        RECT 0.090 279.740 1150.760 281.940 ;
        RECT 0.090 278.580 1150.460 279.740 ;
        RECT 0.090 269.660 1150.760 278.580 ;
        RECT 0.090 268.500 0.700 269.660 ;
        RECT 4.300 268.500 1150.760 269.660 ;
        RECT 0.090 266.300 1150.760 268.500 ;
        RECT 0.090 265.140 1150.460 266.300 ;
        RECT 0.090 259.580 1150.760 265.140 ;
        RECT 0.090 258.420 0.700 259.580 ;
        RECT 4.300 258.420 1150.760 259.580 ;
        RECT 0.090 256.220 1150.760 258.420 ;
        RECT 0.090 255.060 1150.460 256.220 ;
        RECT 0.090 249.500 1150.760 255.060 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 1150.760 249.500 ;
        RECT 0.090 246.140 1150.760 248.340 ;
        RECT 0.090 244.980 1150.460 246.140 ;
        RECT 0.090 236.060 1150.760 244.980 ;
        RECT 0.090 234.900 0.700 236.060 ;
        RECT 4.300 234.900 1150.760 236.060 ;
        RECT 0.090 232.700 1150.760 234.900 ;
        RECT 0.090 231.540 1150.460 232.700 ;
        RECT 0.090 225.980 1150.760 231.540 ;
        RECT 0.090 224.820 0.700 225.980 ;
        RECT 4.300 224.820 1150.760 225.980 ;
        RECT 0.090 222.620 1150.760 224.820 ;
        RECT 0.090 221.460 1150.460 222.620 ;
        RECT 0.090 212.540 1150.760 221.460 ;
        RECT 0.090 211.380 0.700 212.540 ;
        RECT 4.300 211.380 1150.460 212.540 ;
        RECT 0.090 202.460 1150.760 211.380 ;
        RECT 0.090 201.300 0.700 202.460 ;
        RECT 4.300 201.300 1150.760 202.460 ;
        RECT 0.090 199.100 1150.760 201.300 ;
        RECT 0.090 197.940 1150.460 199.100 ;
        RECT 0.090 192.380 1150.760 197.940 ;
        RECT 0.090 191.220 0.700 192.380 ;
        RECT 4.300 191.220 1150.760 192.380 ;
        RECT 0.090 189.020 1150.760 191.220 ;
        RECT 0.090 187.860 1150.460 189.020 ;
        RECT 0.090 178.940 1150.760 187.860 ;
        RECT 0.090 177.780 0.700 178.940 ;
        RECT 4.300 177.780 1150.760 178.940 ;
        RECT 0.090 175.580 1150.760 177.780 ;
        RECT 0.090 174.420 1150.460 175.580 ;
        RECT 0.090 168.860 1150.760 174.420 ;
        RECT 0.090 167.700 0.700 168.860 ;
        RECT 4.300 167.700 1150.760 168.860 ;
        RECT 0.090 165.500 1150.760 167.700 ;
        RECT 0.090 164.340 1150.460 165.500 ;
        RECT 0.090 158.780 1150.760 164.340 ;
        RECT 0.090 157.620 0.700 158.780 ;
        RECT 4.300 157.620 1150.760 158.780 ;
        RECT 0.090 155.420 1150.760 157.620 ;
        RECT 0.090 154.260 1150.460 155.420 ;
        RECT 0.090 145.340 1150.760 154.260 ;
        RECT 0.090 144.180 0.700 145.340 ;
        RECT 4.300 144.180 1150.760 145.340 ;
        RECT 0.090 141.980 1150.760 144.180 ;
        RECT 0.090 140.820 1150.460 141.980 ;
        RECT 0.090 135.260 1150.760 140.820 ;
        RECT 0.090 134.100 0.700 135.260 ;
        RECT 4.300 134.100 1150.760 135.260 ;
        RECT 0.090 131.900 1150.760 134.100 ;
        RECT 0.090 130.740 1150.460 131.900 ;
        RECT 0.090 125.180 1150.760 130.740 ;
        RECT 0.090 124.020 0.700 125.180 ;
        RECT 4.300 124.020 1150.760 125.180 ;
        RECT 0.090 121.820 1150.760 124.020 ;
        RECT 0.090 120.660 1150.460 121.820 ;
        RECT 0.090 111.740 1150.760 120.660 ;
        RECT 0.090 110.580 0.700 111.740 ;
        RECT 4.300 110.580 1150.760 111.740 ;
        RECT 0.090 108.380 1150.760 110.580 ;
        RECT 0.090 107.220 1150.460 108.380 ;
        RECT 0.090 101.660 1150.760 107.220 ;
        RECT 0.090 100.500 0.700 101.660 ;
        RECT 4.300 100.500 1150.760 101.660 ;
        RECT 0.090 98.300 1150.760 100.500 ;
        RECT 0.090 97.140 1150.460 98.300 ;
        RECT 0.090 88.220 1150.760 97.140 ;
        RECT 0.090 87.060 0.700 88.220 ;
        RECT 4.300 87.060 1150.460 88.220 ;
        RECT 0.090 78.140 1150.760 87.060 ;
        RECT 0.090 76.980 0.700 78.140 ;
        RECT 4.300 76.980 1150.760 78.140 ;
        RECT 0.090 74.780 1150.760 76.980 ;
        RECT 0.090 73.620 1150.460 74.780 ;
        RECT 0.090 68.060 1150.760 73.620 ;
        RECT 0.090 66.900 0.700 68.060 ;
        RECT 4.300 66.900 1150.760 68.060 ;
        RECT 0.090 64.700 1150.760 66.900 ;
        RECT 0.090 63.540 1150.460 64.700 ;
        RECT 0.090 54.620 1150.760 63.540 ;
        RECT 0.090 53.460 0.700 54.620 ;
        RECT 4.300 53.460 1150.760 54.620 ;
        RECT 0.090 51.260 1150.760 53.460 ;
        RECT 0.090 50.100 1150.460 51.260 ;
        RECT 0.090 44.540 1150.760 50.100 ;
        RECT 0.090 43.380 0.700 44.540 ;
        RECT 4.300 43.380 1150.760 44.540 ;
        RECT 0.090 41.180 1150.760 43.380 ;
        RECT 0.090 40.020 1150.460 41.180 ;
        RECT 0.090 34.460 1150.760 40.020 ;
        RECT 0.090 33.300 0.700 34.460 ;
        RECT 4.300 33.300 1150.760 34.460 ;
        RECT 0.090 31.100 1150.760 33.300 ;
        RECT 0.090 29.940 1150.460 31.100 ;
        RECT 0.090 21.020 1150.760 29.940 ;
        RECT 0.090 19.860 0.700 21.020 ;
        RECT 4.300 19.860 1150.760 21.020 ;
        RECT 0.090 17.660 1150.760 19.860 ;
        RECT 0.090 16.500 1150.460 17.660 ;
        RECT 0.090 10.940 1150.760 16.500 ;
        RECT 0.090 9.780 0.700 10.940 ;
        RECT 4.300 9.780 1150.760 10.940 ;
        RECT 0.090 9.100 1150.760 9.780 ;
      LAYER Metal4 ;
        RECT 61.740 17.450 98.740 1154.630 ;
        RECT 100.940 17.450 175.540 1154.630 ;
        RECT 177.740 17.450 252.340 1154.630 ;
        RECT 254.540 17.450 329.140 1154.630 ;
        RECT 331.340 17.450 405.940 1154.630 ;
        RECT 408.140 17.450 482.740 1154.630 ;
        RECT 484.940 17.450 559.540 1154.630 ;
        RECT 561.740 17.450 636.340 1154.630 ;
        RECT 638.540 17.450 713.140 1154.630 ;
        RECT 715.340 17.450 789.940 1154.630 ;
        RECT 792.140 17.450 866.740 1154.630 ;
        RECT 868.940 17.450 943.540 1154.630 ;
        RECT 945.740 17.450 1020.340 1154.630 ;
        RECT 1022.540 17.450 1097.140 1154.630 ;
        RECT 1099.340 17.450 1139.460 1154.630 ;
  END
END aes_core
END LIBRARY

