magic
tech gf180mcuC
magscale 1 5
timestamp 1669631042
<< obsm1 >>
rect 672 855 114800 115737
<< metal2 >>
rect 0 116868 56 117168
rect 1344 116868 1400 117168
rect 2352 116868 2408 117168
rect 3360 116868 3416 117168
rect 4704 116868 4760 117168
rect 5712 116868 5768 117168
rect 7056 116868 7112 117168
rect 8064 116868 8120 117168
rect 9072 116868 9128 117168
rect 10416 116868 10472 117168
rect 11424 116868 11480 117168
rect 12432 116868 12488 117168
rect 13776 116868 13832 117168
rect 14784 116868 14840 117168
rect 15792 116868 15848 117168
rect 17136 116868 17192 117168
rect 18144 116868 18200 117168
rect 19488 116868 19544 117168
rect 20496 116868 20552 117168
rect 21504 116868 21560 117168
rect 22848 116868 22904 117168
rect 23856 116868 23912 117168
rect 24864 116868 24920 117168
rect 26208 116868 26264 117168
rect 27216 116868 27272 117168
rect 28224 116868 28280 117168
rect 29568 116868 29624 117168
rect 30576 116868 30632 117168
rect 31920 116868 31976 117168
rect 32928 116868 32984 117168
rect 33936 116868 33992 117168
rect 35280 116868 35336 117168
rect 36288 116868 36344 117168
rect 37296 116868 37352 117168
rect 38640 116868 38696 117168
rect 39648 116868 39704 117168
rect 40656 116868 40712 117168
rect 42000 116868 42056 117168
rect 43008 116868 43064 117168
rect 44352 116868 44408 117168
rect 45360 116868 45416 117168
rect 46368 116868 46424 117168
rect 47712 116868 47768 117168
rect 48720 116868 48776 117168
rect 49728 116868 49784 117168
rect 51072 116868 51128 117168
rect 52080 116868 52136 117168
rect 53088 116868 53144 117168
rect 54432 116868 54488 117168
rect 55440 116868 55496 117168
rect 56784 116868 56840 117168
rect 57792 116868 57848 117168
rect 58800 116868 58856 117168
rect 60144 116868 60200 117168
rect 61152 116868 61208 117168
rect 62160 116868 62216 117168
rect 63504 116868 63560 117168
rect 64512 116868 64568 117168
rect 65520 116868 65576 117168
rect 66864 116868 66920 117168
rect 67872 116868 67928 117168
rect 69216 116868 69272 117168
rect 70224 116868 70280 117168
rect 71232 116868 71288 117168
rect 72576 116868 72632 117168
rect 73584 116868 73640 117168
rect 74592 116868 74648 117168
rect 75936 116868 75992 117168
rect 76944 116868 77000 117168
rect 77952 116868 78008 117168
rect 79296 116868 79352 117168
rect 80304 116868 80360 117168
rect 81648 116868 81704 117168
rect 82656 116868 82712 117168
rect 83664 116868 83720 117168
rect 85008 116868 85064 117168
rect 86016 116868 86072 117168
rect 87024 116868 87080 117168
rect 88368 116868 88424 117168
rect 89376 116868 89432 117168
rect 90384 116868 90440 117168
rect 91728 116868 91784 117168
rect 92736 116868 92792 117168
rect 94080 116868 94136 117168
rect 95088 116868 95144 117168
rect 96096 116868 96152 117168
rect 97440 116868 97496 117168
rect 98448 116868 98504 117168
rect 99456 116868 99512 117168
rect 100800 116868 100856 117168
rect 101808 116868 101864 117168
rect 102816 116868 102872 117168
rect 104160 116868 104216 117168
rect 105168 116868 105224 117168
rect 106512 116868 106568 117168
rect 107520 116868 107576 117168
rect 108528 116868 108584 117168
rect 109872 116868 109928 117168
rect 110880 116868 110936 117168
rect 111888 116868 111944 117168
rect 113232 116868 113288 117168
rect 114240 116868 114296 117168
rect 115248 116868 115304 117168
rect 0 100 56 400
rect 1008 100 1064 400
rect 2016 100 2072 400
rect 3360 100 3416 400
rect 4368 100 4424 400
rect 5376 100 5432 400
rect 6720 100 6776 400
rect 7728 100 7784 400
rect 8736 100 8792 400
rect 10080 100 10136 400
rect 11088 100 11144 400
rect 12432 100 12488 400
rect 13440 100 13496 400
rect 14448 100 14504 400
rect 15792 100 15848 400
rect 16800 100 16856 400
rect 17808 100 17864 400
rect 19152 100 19208 400
rect 20160 100 20216 400
rect 21168 100 21224 400
rect 22512 100 22568 400
rect 23520 100 23576 400
rect 24864 100 24920 400
rect 25872 100 25928 400
rect 26880 100 26936 400
rect 28224 100 28280 400
rect 29232 100 29288 400
rect 30240 100 30296 400
rect 31584 100 31640 400
rect 32592 100 32648 400
rect 33600 100 33656 400
rect 34944 100 35000 400
rect 35952 100 36008 400
rect 37296 100 37352 400
rect 38304 100 38360 400
rect 39312 100 39368 400
rect 40656 100 40712 400
rect 41664 100 41720 400
rect 42672 100 42728 400
rect 44016 100 44072 400
rect 45024 100 45080 400
rect 46032 100 46088 400
rect 47376 100 47432 400
rect 48384 100 48440 400
rect 49728 100 49784 400
rect 50736 100 50792 400
rect 51744 100 51800 400
rect 53088 100 53144 400
rect 54096 100 54152 400
rect 55104 100 55160 400
rect 56448 100 56504 400
rect 57456 100 57512 400
rect 58464 100 58520 400
rect 59808 100 59864 400
rect 60816 100 60872 400
rect 62160 100 62216 400
rect 63168 100 63224 400
rect 64176 100 64232 400
rect 65520 100 65576 400
rect 66528 100 66584 400
rect 67536 100 67592 400
rect 68880 100 68936 400
rect 69888 100 69944 400
rect 70896 100 70952 400
rect 72240 100 72296 400
rect 73248 100 73304 400
rect 74592 100 74648 400
rect 75600 100 75656 400
rect 76608 100 76664 400
rect 77952 100 78008 400
rect 78960 100 79016 400
rect 79968 100 80024 400
rect 81312 100 81368 400
rect 82320 100 82376 400
rect 83328 100 83384 400
rect 84672 100 84728 400
rect 85680 100 85736 400
rect 87024 100 87080 400
rect 88032 100 88088 400
rect 89040 100 89096 400
rect 90384 100 90440 400
rect 91392 100 91448 400
rect 92400 100 92456 400
rect 93744 100 93800 400
rect 94752 100 94808 400
rect 95760 100 95816 400
rect 97104 100 97160 400
rect 98112 100 98168 400
rect 99456 100 99512 400
rect 100464 100 100520 400
rect 101472 100 101528 400
rect 102816 100 102872 400
rect 103824 100 103880 400
rect 104832 100 104888 400
rect 106176 100 106232 400
rect 107184 100 107240 400
rect 108192 100 108248 400
rect 109536 100 109592 400
rect 110544 100 110600 400
rect 111888 100 111944 400
rect 112896 100 112952 400
rect 113904 100 113960 400
rect 115248 100 115304 400
<< obsm2 >>
rect 86 116838 1314 116914
rect 1430 116838 2322 116914
rect 2438 116838 3330 116914
rect 3446 116838 4674 116914
rect 4790 116838 5682 116914
rect 5798 116838 7026 116914
rect 7142 116838 8034 116914
rect 8150 116838 9042 116914
rect 9158 116838 10386 116914
rect 10502 116838 11394 116914
rect 11510 116838 12402 116914
rect 12518 116838 13746 116914
rect 13862 116838 14754 116914
rect 14870 116838 15762 116914
rect 15878 116838 17106 116914
rect 17222 116838 18114 116914
rect 18230 116838 19458 116914
rect 19574 116838 20466 116914
rect 20582 116838 21474 116914
rect 21590 116838 22818 116914
rect 22934 116838 23826 116914
rect 23942 116838 24834 116914
rect 24950 116838 26178 116914
rect 26294 116838 27186 116914
rect 27302 116838 28194 116914
rect 28310 116838 29538 116914
rect 29654 116838 30546 116914
rect 30662 116838 31890 116914
rect 32006 116838 32898 116914
rect 33014 116838 33906 116914
rect 34022 116838 35250 116914
rect 35366 116838 36258 116914
rect 36374 116838 37266 116914
rect 37382 116838 38610 116914
rect 38726 116838 39618 116914
rect 39734 116838 40626 116914
rect 40742 116838 41970 116914
rect 42086 116838 42978 116914
rect 43094 116838 44322 116914
rect 44438 116838 45330 116914
rect 45446 116838 46338 116914
rect 46454 116838 47682 116914
rect 47798 116838 48690 116914
rect 48806 116838 49698 116914
rect 49814 116838 51042 116914
rect 51158 116838 52050 116914
rect 52166 116838 53058 116914
rect 53174 116838 54402 116914
rect 54518 116838 55410 116914
rect 55526 116838 56754 116914
rect 56870 116838 57762 116914
rect 57878 116838 58770 116914
rect 58886 116838 60114 116914
rect 60230 116838 61122 116914
rect 61238 116838 62130 116914
rect 62246 116838 63474 116914
rect 63590 116838 64482 116914
rect 64598 116838 65490 116914
rect 65606 116838 66834 116914
rect 66950 116838 67842 116914
rect 67958 116838 69186 116914
rect 69302 116838 70194 116914
rect 70310 116838 71202 116914
rect 71318 116838 72546 116914
rect 72662 116838 73554 116914
rect 73670 116838 74562 116914
rect 74678 116838 75906 116914
rect 76022 116838 76914 116914
rect 77030 116838 77922 116914
rect 78038 116838 79266 116914
rect 79382 116838 80274 116914
rect 80390 116838 81618 116914
rect 81734 116838 82626 116914
rect 82742 116838 83634 116914
rect 83750 116838 84978 116914
rect 85094 116838 85986 116914
rect 86102 116838 86994 116914
rect 87110 116838 88338 116914
rect 88454 116838 89346 116914
rect 89462 116838 90354 116914
rect 90470 116838 91698 116914
rect 91814 116838 92706 116914
rect 92822 116838 94050 116914
rect 94166 116838 95058 116914
rect 95174 116838 96066 116914
rect 96182 116838 97410 116914
rect 97526 116838 98418 116914
rect 98534 116838 99426 116914
rect 99542 116838 100770 116914
rect 100886 116838 101778 116914
rect 101894 116838 102786 116914
rect 102902 116838 104130 116914
rect 104246 116838 105138 116914
rect 105254 116838 106482 116914
rect 106598 116838 107490 116914
rect 107606 116838 108498 116914
rect 108614 116838 109842 116914
rect 109958 116838 110850 116914
rect 110966 116838 111858 116914
rect 111974 116838 113202 116914
rect 113318 116838 114210 116914
rect 114326 116838 114674 116914
rect 14 430 114674 116838
rect 86 400 978 430
rect 1094 400 1986 430
rect 2102 400 3330 430
rect 3446 400 4338 430
rect 4454 400 5346 430
rect 5462 400 6690 430
rect 6806 400 7698 430
rect 7814 400 8706 430
rect 8822 400 10050 430
rect 10166 400 11058 430
rect 11174 400 12402 430
rect 12518 400 13410 430
rect 13526 400 14418 430
rect 14534 400 15762 430
rect 15878 400 16770 430
rect 16886 400 17778 430
rect 17894 400 19122 430
rect 19238 400 20130 430
rect 20246 400 21138 430
rect 21254 400 22482 430
rect 22598 400 23490 430
rect 23606 400 24834 430
rect 24950 400 25842 430
rect 25958 400 26850 430
rect 26966 400 28194 430
rect 28310 400 29202 430
rect 29318 400 30210 430
rect 30326 400 31554 430
rect 31670 400 32562 430
rect 32678 400 33570 430
rect 33686 400 34914 430
rect 35030 400 35922 430
rect 36038 400 37266 430
rect 37382 400 38274 430
rect 38390 400 39282 430
rect 39398 400 40626 430
rect 40742 400 41634 430
rect 41750 400 42642 430
rect 42758 400 43986 430
rect 44102 400 44994 430
rect 45110 400 46002 430
rect 46118 400 47346 430
rect 47462 400 48354 430
rect 48470 400 49698 430
rect 49814 400 50706 430
rect 50822 400 51714 430
rect 51830 400 53058 430
rect 53174 400 54066 430
rect 54182 400 55074 430
rect 55190 400 56418 430
rect 56534 400 57426 430
rect 57542 400 58434 430
rect 58550 400 59778 430
rect 59894 400 60786 430
rect 60902 400 62130 430
rect 62246 400 63138 430
rect 63254 400 64146 430
rect 64262 400 65490 430
rect 65606 400 66498 430
rect 66614 400 67506 430
rect 67622 400 68850 430
rect 68966 400 69858 430
rect 69974 400 70866 430
rect 70982 400 72210 430
rect 72326 400 73218 430
rect 73334 400 74562 430
rect 74678 400 75570 430
rect 75686 400 76578 430
rect 76694 400 77922 430
rect 78038 400 78930 430
rect 79046 400 79938 430
rect 80054 400 81282 430
rect 81398 400 82290 430
rect 82406 400 83298 430
rect 83414 400 84642 430
rect 84758 400 85650 430
rect 85766 400 86994 430
rect 87110 400 88002 430
rect 88118 400 89010 430
rect 89126 400 90354 430
rect 90470 400 91362 430
rect 91478 400 92370 430
rect 92486 400 93714 430
rect 93830 400 94722 430
rect 94838 400 95730 430
rect 95846 400 97074 430
rect 97190 400 98082 430
rect 98198 400 99426 430
rect 99542 400 100434 430
rect 100550 400 101442 430
rect 101558 400 102786 430
rect 102902 400 103794 430
rect 103910 400 104802 430
rect 104918 400 106146 430
rect 106262 400 107154 430
rect 107270 400 108162 430
rect 108278 400 109506 430
rect 109622 400 110514 430
rect 110630 400 111858 430
rect 111974 400 112866 430
rect 112982 400 113874 430
rect 113990 400 114674 430
<< metal3 >>
rect 100 116256 400 116312
rect 115076 115920 115376 115976
rect 100 115248 400 115304
rect 115076 114912 115376 114968
rect 100 113904 400 113960
rect 115076 113568 115376 113624
rect 100 112896 400 112952
rect 115076 112560 115376 112616
rect 100 111888 400 111944
rect 115076 111552 115376 111608
rect 100 110544 400 110600
rect 115076 110208 115376 110264
rect 100 109536 400 109592
rect 115076 109200 115376 109256
rect 100 108192 400 108248
rect 115076 108192 115376 108248
rect 100 107184 400 107240
rect 115076 106848 115376 106904
rect 100 106176 400 106232
rect 115076 105840 115376 105896
rect 100 104832 400 104888
rect 115076 104496 115376 104552
rect 100 103824 400 103880
rect 115076 103488 115376 103544
rect 100 102816 400 102872
rect 115076 102480 115376 102536
rect 100 101472 400 101528
rect 115076 101136 115376 101192
rect 100 100464 400 100520
rect 115076 100128 115376 100184
rect 100 99456 400 99512
rect 115076 99120 115376 99176
rect 100 98112 400 98168
rect 115076 97776 115376 97832
rect 100 97104 400 97160
rect 115076 96768 115376 96824
rect 100 95760 400 95816
rect 115076 95760 115376 95816
rect 100 94752 400 94808
rect 115076 94416 115376 94472
rect 100 93744 400 93800
rect 115076 93408 115376 93464
rect 100 92400 400 92456
rect 115076 92064 115376 92120
rect 100 91392 400 91448
rect 115076 91056 115376 91112
rect 100 90384 400 90440
rect 115076 90048 115376 90104
rect 100 89040 400 89096
rect 115076 88704 115376 88760
rect 100 88032 400 88088
rect 115076 87696 115376 87752
rect 100 87024 400 87080
rect 115076 86688 115376 86744
rect 100 85680 400 85736
rect 115076 85344 115376 85400
rect 100 84672 400 84728
rect 115076 84336 115376 84392
rect 100 83328 400 83384
rect 115076 83328 115376 83384
rect 100 82320 400 82376
rect 115076 81984 115376 82040
rect 100 81312 400 81368
rect 115076 80976 115376 81032
rect 100 79968 400 80024
rect 115076 79632 115376 79688
rect 100 78960 400 79016
rect 115076 78624 115376 78680
rect 100 77952 400 78008
rect 115076 77616 115376 77672
rect 100 76608 400 76664
rect 115076 76272 115376 76328
rect 100 75600 400 75656
rect 115076 75264 115376 75320
rect 100 74592 400 74648
rect 115076 74256 115376 74312
rect 100 73248 400 73304
rect 115076 72912 115376 72968
rect 100 72240 400 72296
rect 115076 71904 115376 71960
rect 100 70896 400 70952
rect 115076 70896 115376 70952
rect 100 69888 400 69944
rect 115076 69552 115376 69608
rect 100 68880 400 68936
rect 115076 68544 115376 68600
rect 100 67536 400 67592
rect 115076 67200 115376 67256
rect 100 66528 400 66584
rect 115076 66192 115376 66248
rect 100 65520 400 65576
rect 115076 65184 115376 65240
rect 100 64176 400 64232
rect 115076 63840 115376 63896
rect 100 63168 400 63224
rect 115076 62832 115376 62888
rect 100 62160 400 62216
rect 115076 61824 115376 61880
rect 100 60816 400 60872
rect 115076 60480 115376 60536
rect 100 59808 400 59864
rect 115076 59472 115376 59528
rect 100 58464 400 58520
rect 115076 58464 115376 58520
rect 100 57456 400 57512
rect 115076 57120 115376 57176
rect 100 56448 400 56504
rect 115076 56112 115376 56168
rect 100 55104 400 55160
rect 115076 54768 115376 54824
rect 100 54096 400 54152
rect 115076 53760 115376 53816
rect 100 53088 400 53144
rect 115076 52752 115376 52808
rect 100 51744 400 51800
rect 115076 51408 115376 51464
rect 100 50736 400 50792
rect 115076 50400 115376 50456
rect 100 49728 400 49784
rect 115076 49392 115376 49448
rect 100 48384 400 48440
rect 115076 48048 115376 48104
rect 100 47376 400 47432
rect 115076 47040 115376 47096
rect 100 46032 400 46088
rect 115076 46032 115376 46088
rect 100 45024 400 45080
rect 115076 44688 115376 44744
rect 100 44016 400 44072
rect 115076 43680 115376 43736
rect 100 42672 400 42728
rect 115076 42336 115376 42392
rect 100 41664 400 41720
rect 115076 41328 115376 41384
rect 100 40656 400 40712
rect 115076 40320 115376 40376
rect 100 39312 400 39368
rect 115076 38976 115376 39032
rect 100 38304 400 38360
rect 115076 37968 115376 38024
rect 100 37296 400 37352
rect 115076 36960 115376 37016
rect 100 35952 400 36008
rect 115076 35616 115376 35672
rect 100 34944 400 35000
rect 115076 34608 115376 34664
rect 100 33600 400 33656
rect 115076 33600 115376 33656
rect 100 32592 400 32648
rect 115076 32256 115376 32312
rect 100 31584 400 31640
rect 115076 31248 115376 31304
rect 100 30240 400 30296
rect 115076 29904 115376 29960
rect 100 29232 400 29288
rect 115076 28896 115376 28952
rect 100 28224 400 28280
rect 115076 27888 115376 27944
rect 100 26880 400 26936
rect 115076 26544 115376 26600
rect 100 25872 400 25928
rect 115076 25536 115376 25592
rect 100 24864 400 24920
rect 115076 24528 115376 24584
rect 100 23520 400 23576
rect 115076 23184 115376 23240
rect 100 22512 400 22568
rect 115076 22176 115376 22232
rect 100 21168 400 21224
rect 115076 21168 115376 21224
rect 100 20160 400 20216
rect 115076 19824 115376 19880
rect 100 19152 400 19208
rect 115076 18816 115376 18872
rect 100 17808 400 17864
rect 115076 17472 115376 17528
rect 100 16800 400 16856
rect 115076 16464 115376 16520
rect 100 15792 400 15848
rect 115076 15456 115376 15512
rect 100 14448 400 14504
rect 115076 14112 115376 14168
rect 100 13440 400 13496
rect 115076 13104 115376 13160
rect 100 12432 400 12488
rect 115076 12096 115376 12152
rect 100 11088 400 11144
rect 115076 10752 115376 10808
rect 100 10080 400 10136
rect 115076 9744 115376 9800
rect 100 8736 400 8792
rect 115076 8736 115376 8792
rect 100 7728 400 7784
rect 115076 7392 115376 7448
rect 100 6720 400 6776
rect 115076 6384 115376 6440
rect 100 5376 400 5432
rect 115076 5040 115376 5096
rect 100 4368 400 4424
rect 115076 4032 115376 4088
rect 100 3360 400 3416
rect 115076 3024 115376 3080
rect 100 2016 400 2072
rect 115076 1680 115376 1736
rect 100 1008 400 1064
rect 115076 672 115376 728
<< obsm3 >>
rect 9 115334 115076 115738
rect 9 115218 70 115334
rect 430 115218 115076 115334
rect 9 114998 115076 115218
rect 9 114882 115046 114998
rect 9 113990 115076 114882
rect 9 113874 70 113990
rect 430 113874 115076 113990
rect 9 113654 115076 113874
rect 9 113538 115046 113654
rect 9 112982 115076 113538
rect 9 112866 70 112982
rect 430 112866 115076 112982
rect 9 112646 115076 112866
rect 9 112530 115046 112646
rect 9 111974 115076 112530
rect 9 111858 70 111974
rect 430 111858 115076 111974
rect 9 111638 115076 111858
rect 9 111522 115046 111638
rect 9 110630 115076 111522
rect 9 110514 70 110630
rect 430 110514 115076 110630
rect 9 110294 115076 110514
rect 9 110178 115046 110294
rect 9 109622 115076 110178
rect 9 109506 70 109622
rect 430 109506 115076 109622
rect 9 109286 115076 109506
rect 9 109170 115046 109286
rect 9 108278 115076 109170
rect 9 108162 70 108278
rect 430 108162 115046 108278
rect 9 107270 115076 108162
rect 9 107154 70 107270
rect 430 107154 115076 107270
rect 9 106934 115076 107154
rect 9 106818 115046 106934
rect 9 106262 115076 106818
rect 9 106146 70 106262
rect 430 106146 115076 106262
rect 9 105926 115076 106146
rect 9 105810 115046 105926
rect 9 104918 115076 105810
rect 9 104802 70 104918
rect 430 104802 115076 104918
rect 9 104582 115076 104802
rect 9 104466 115046 104582
rect 9 103910 115076 104466
rect 9 103794 70 103910
rect 430 103794 115076 103910
rect 9 103574 115076 103794
rect 9 103458 115046 103574
rect 9 102902 115076 103458
rect 9 102786 70 102902
rect 430 102786 115076 102902
rect 9 102566 115076 102786
rect 9 102450 115046 102566
rect 9 101558 115076 102450
rect 9 101442 70 101558
rect 430 101442 115076 101558
rect 9 101222 115076 101442
rect 9 101106 115046 101222
rect 9 100550 115076 101106
rect 9 100434 70 100550
rect 430 100434 115076 100550
rect 9 100214 115076 100434
rect 9 100098 115046 100214
rect 9 99542 115076 100098
rect 9 99426 70 99542
rect 430 99426 115076 99542
rect 9 99206 115076 99426
rect 9 99090 115046 99206
rect 9 98198 115076 99090
rect 9 98082 70 98198
rect 430 98082 115076 98198
rect 9 97862 115076 98082
rect 9 97746 115046 97862
rect 9 97190 115076 97746
rect 9 97074 70 97190
rect 430 97074 115076 97190
rect 9 96854 115076 97074
rect 9 96738 115046 96854
rect 9 95846 115076 96738
rect 9 95730 70 95846
rect 430 95730 115046 95846
rect 9 94838 115076 95730
rect 9 94722 70 94838
rect 430 94722 115076 94838
rect 9 94502 115076 94722
rect 9 94386 115046 94502
rect 9 93830 115076 94386
rect 9 93714 70 93830
rect 430 93714 115076 93830
rect 9 93494 115076 93714
rect 9 93378 115046 93494
rect 9 92486 115076 93378
rect 9 92370 70 92486
rect 430 92370 115076 92486
rect 9 92150 115076 92370
rect 9 92034 115046 92150
rect 9 91478 115076 92034
rect 9 91362 70 91478
rect 430 91362 115076 91478
rect 9 91142 115076 91362
rect 9 91026 115046 91142
rect 9 90470 115076 91026
rect 9 90354 70 90470
rect 430 90354 115076 90470
rect 9 90134 115076 90354
rect 9 90018 115046 90134
rect 9 89126 115076 90018
rect 9 89010 70 89126
rect 430 89010 115076 89126
rect 9 88790 115076 89010
rect 9 88674 115046 88790
rect 9 88118 115076 88674
rect 9 88002 70 88118
rect 430 88002 115076 88118
rect 9 87782 115076 88002
rect 9 87666 115046 87782
rect 9 87110 115076 87666
rect 9 86994 70 87110
rect 430 86994 115076 87110
rect 9 86774 115076 86994
rect 9 86658 115046 86774
rect 9 85766 115076 86658
rect 9 85650 70 85766
rect 430 85650 115076 85766
rect 9 85430 115076 85650
rect 9 85314 115046 85430
rect 9 84758 115076 85314
rect 9 84642 70 84758
rect 430 84642 115076 84758
rect 9 84422 115076 84642
rect 9 84306 115046 84422
rect 9 83414 115076 84306
rect 9 83298 70 83414
rect 430 83298 115046 83414
rect 9 82406 115076 83298
rect 9 82290 70 82406
rect 430 82290 115076 82406
rect 9 82070 115076 82290
rect 9 81954 115046 82070
rect 9 81398 115076 81954
rect 9 81282 70 81398
rect 430 81282 115076 81398
rect 9 81062 115076 81282
rect 9 80946 115046 81062
rect 9 80054 115076 80946
rect 9 79938 70 80054
rect 430 79938 115076 80054
rect 9 79718 115076 79938
rect 9 79602 115046 79718
rect 9 79046 115076 79602
rect 9 78930 70 79046
rect 430 78930 115076 79046
rect 9 78710 115076 78930
rect 9 78594 115046 78710
rect 9 78038 115076 78594
rect 9 77922 70 78038
rect 430 77922 115076 78038
rect 9 77702 115076 77922
rect 9 77586 115046 77702
rect 9 76694 115076 77586
rect 9 76578 70 76694
rect 430 76578 115076 76694
rect 9 76358 115076 76578
rect 9 76242 115046 76358
rect 9 75686 115076 76242
rect 9 75570 70 75686
rect 430 75570 115076 75686
rect 9 75350 115076 75570
rect 9 75234 115046 75350
rect 9 74678 115076 75234
rect 9 74562 70 74678
rect 430 74562 115076 74678
rect 9 74342 115076 74562
rect 9 74226 115046 74342
rect 9 73334 115076 74226
rect 9 73218 70 73334
rect 430 73218 115076 73334
rect 9 72998 115076 73218
rect 9 72882 115046 72998
rect 9 72326 115076 72882
rect 9 72210 70 72326
rect 430 72210 115076 72326
rect 9 71990 115076 72210
rect 9 71874 115046 71990
rect 9 70982 115076 71874
rect 9 70866 70 70982
rect 430 70866 115046 70982
rect 9 69974 115076 70866
rect 9 69858 70 69974
rect 430 69858 115076 69974
rect 9 69638 115076 69858
rect 9 69522 115046 69638
rect 9 68966 115076 69522
rect 9 68850 70 68966
rect 430 68850 115076 68966
rect 9 68630 115076 68850
rect 9 68514 115046 68630
rect 9 67622 115076 68514
rect 9 67506 70 67622
rect 430 67506 115076 67622
rect 9 67286 115076 67506
rect 9 67170 115046 67286
rect 9 66614 115076 67170
rect 9 66498 70 66614
rect 430 66498 115076 66614
rect 9 66278 115076 66498
rect 9 66162 115046 66278
rect 9 65606 115076 66162
rect 9 65490 70 65606
rect 430 65490 115076 65606
rect 9 65270 115076 65490
rect 9 65154 115046 65270
rect 9 64262 115076 65154
rect 9 64146 70 64262
rect 430 64146 115076 64262
rect 9 63926 115076 64146
rect 9 63810 115046 63926
rect 9 63254 115076 63810
rect 9 63138 70 63254
rect 430 63138 115076 63254
rect 9 62918 115076 63138
rect 9 62802 115046 62918
rect 9 62246 115076 62802
rect 9 62130 70 62246
rect 430 62130 115076 62246
rect 9 61910 115076 62130
rect 9 61794 115046 61910
rect 9 60902 115076 61794
rect 9 60786 70 60902
rect 430 60786 115076 60902
rect 9 60566 115076 60786
rect 9 60450 115046 60566
rect 9 59894 115076 60450
rect 9 59778 70 59894
rect 430 59778 115076 59894
rect 9 59558 115076 59778
rect 9 59442 115046 59558
rect 9 58550 115076 59442
rect 9 58434 70 58550
rect 430 58434 115046 58550
rect 9 57542 115076 58434
rect 9 57426 70 57542
rect 430 57426 115076 57542
rect 9 57206 115076 57426
rect 9 57090 115046 57206
rect 9 56534 115076 57090
rect 9 56418 70 56534
rect 430 56418 115076 56534
rect 9 56198 115076 56418
rect 9 56082 115046 56198
rect 9 55190 115076 56082
rect 9 55074 70 55190
rect 430 55074 115076 55190
rect 9 54854 115076 55074
rect 9 54738 115046 54854
rect 9 54182 115076 54738
rect 9 54066 70 54182
rect 430 54066 115076 54182
rect 9 53846 115076 54066
rect 9 53730 115046 53846
rect 9 53174 115076 53730
rect 9 53058 70 53174
rect 430 53058 115076 53174
rect 9 52838 115076 53058
rect 9 52722 115046 52838
rect 9 51830 115076 52722
rect 9 51714 70 51830
rect 430 51714 115076 51830
rect 9 51494 115076 51714
rect 9 51378 115046 51494
rect 9 50822 115076 51378
rect 9 50706 70 50822
rect 430 50706 115076 50822
rect 9 50486 115076 50706
rect 9 50370 115046 50486
rect 9 49814 115076 50370
rect 9 49698 70 49814
rect 430 49698 115076 49814
rect 9 49478 115076 49698
rect 9 49362 115046 49478
rect 9 48470 115076 49362
rect 9 48354 70 48470
rect 430 48354 115076 48470
rect 9 48134 115076 48354
rect 9 48018 115046 48134
rect 9 47462 115076 48018
rect 9 47346 70 47462
rect 430 47346 115076 47462
rect 9 47126 115076 47346
rect 9 47010 115046 47126
rect 9 46118 115076 47010
rect 9 46002 70 46118
rect 430 46002 115046 46118
rect 9 45110 115076 46002
rect 9 44994 70 45110
rect 430 44994 115076 45110
rect 9 44774 115076 44994
rect 9 44658 115046 44774
rect 9 44102 115076 44658
rect 9 43986 70 44102
rect 430 43986 115076 44102
rect 9 43766 115076 43986
rect 9 43650 115046 43766
rect 9 42758 115076 43650
rect 9 42642 70 42758
rect 430 42642 115076 42758
rect 9 42422 115076 42642
rect 9 42306 115046 42422
rect 9 41750 115076 42306
rect 9 41634 70 41750
rect 430 41634 115076 41750
rect 9 41414 115076 41634
rect 9 41298 115046 41414
rect 9 40742 115076 41298
rect 9 40626 70 40742
rect 430 40626 115076 40742
rect 9 40406 115076 40626
rect 9 40290 115046 40406
rect 9 39398 115076 40290
rect 9 39282 70 39398
rect 430 39282 115076 39398
rect 9 39062 115076 39282
rect 9 38946 115046 39062
rect 9 38390 115076 38946
rect 9 38274 70 38390
rect 430 38274 115076 38390
rect 9 38054 115076 38274
rect 9 37938 115046 38054
rect 9 37382 115076 37938
rect 9 37266 70 37382
rect 430 37266 115076 37382
rect 9 37046 115076 37266
rect 9 36930 115046 37046
rect 9 36038 115076 36930
rect 9 35922 70 36038
rect 430 35922 115076 36038
rect 9 35702 115076 35922
rect 9 35586 115046 35702
rect 9 35030 115076 35586
rect 9 34914 70 35030
rect 430 34914 115076 35030
rect 9 34694 115076 34914
rect 9 34578 115046 34694
rect 9 33686 115076 34578
rect 9 33570 70 33686
rect 430 33570 115046 33686
rect 9 32678 115076 33570
rect 9 32562 70 32678
rect 430 32562 115076 32678
rect 9 32342 115076 32562
rect 9 32226 115046 32342
rect 9 31670 115076 32226
rect 9 31554 70 31670
rect 430 31554 115076 31670
rect 9 31334 115076 31554
rect 9 31218 115046 31334
rect 9 30326 115076 31218
rect 9 30210 70 30326
rect 430 30210 115076 30326
rect 9 29990 115076 30210
rect 9 29874 115046 29990
rect 9 29318 115076 29874
rect 9 29202 70 29318
rect 430 29202 115076 29318
rect 9 28982 115076 29202
rect 9 28866 115046 28982
rect 9 28310 115076 28866
rect 9 28194 70 28310
rect 430 28194 115076 28310
rect 9 27974 115076 28194
rect 9 27858 115046 27974
rect 9 26966 115076 27858
rect 9 26850 70 26966
rect 430 26850 115076 26966
rect 9 26630 115076 26850
rect 9 26514 115046 26630
rect 9 25958 115076 26514
rect 9 25842 70 25958
rect 430 25842 115076 25958
rect 9 25622 115076 25842
rect 9 25506 115046 25622
rect 9 24950 115076 25506
rect 9 24834 70 24950
rect 430 24834 115076 24950
rect 9 24614 115076 24834
rect 9 24498 115046 24614
rect 9 23606 115076 24498
rect 9 23490 70 23606
rect 430 23490 115076 23606
rect 9 23270 115076 23490
rect 9 23154 115046 23270
rect 9 22598 115076 23154
rect 9 22482 70 22598
rect 430 22482 115076 22598
rect 9 22262 115076 22482
rect 9 22146 115046 22262
rect 9 21254 115076 22146
rect 9 21138 70 21254
rect 430 21138 115046 21254
rect 9 20246 115076 21138
rect 9 20130 70 20246
rect 430 20130 115076 20246
rect 9 19910 115076 20130
rect 9 19794 115046 19910
rect 9 19238 115076 19794
rect 9 19122 70 19238
rect 430 19122 115076 19238
rect 9 18902 115076 19122
rect 9 18786 115046 18902
rect 9 17894 115076 18786
rect 9 17778 70 17894
rect 430 17778 115076 17894
rect 9 17558 115076 17778
rect 9 17442 115046 17558
rect 9 16886 115076 17442
rect 9 16770 70 16886
rect 430 16770 115076 16886
rect 9 16550 115076 16770
rect 9 16434 115046 16550
rect 9 15878 115076 16434
rect 9 15762 70 15878
rect 430 15762 115076 15878
rect 9 15542 115076 15762
rect 9 15426 115046 15542
rect 9 14534 115076 15426
rect 9 14418 70 14534
rect 430 14418 115076 14534
rect 9 14198 115076 14418
rect 9 14082 115046 14198
rect 9 13526 115076 14082
rect 9 13410 70 13526
rect 430 13410 115076 13526
rect 9 13190 115076 13410
rect 9 13074 115046 13190
rect 9 12518 115076 13074
rect 9 12402 70 12518
rect 430 12402 115076 12518
rect 9 12182 115076 12402
rect 9 12066 115046 12182
rect 9 11174 115076 12066
rect 9 11058 70 11174
rect 430 11058 115076 11174
rect 9 10838 115076 11058
rect 9 10722 115046 10838
rect 9 10166 115076 10722
rect 9 10050 70 10166
rect 430 10050 115076 10166
rect 9 9830 115076 10050
rect 9 9714 115046 9830
rect 9 8822 115076 9714
rect 9 8706 70 8822
rect 430 8706 115046 8822
rect 9 7814 115076 8706
rect 9 7698 70 7814
rect 430 7698 115076 7814
rect 9 7478 115076 7698
rect 9 7362 115046 7478
rect 9 6806 115076 7362
rect 9 6690 70 6806
rect 430 6690 115076 6806
rect 9 6470 115076 6690
rect 9 6354 115046 6470
rect 9 5462 115076 6354
rect 9 5346 70 5462
rect 430 5346 115076 5462
rect 9 5126 115076 5346
rect 9 5010 115046 5126
rect 9 4454 115076 5010
rect 9 4338 70 4454
rect 430 4338 115076 4454
rect 9 4118 115076 4338
rect 9 4002 115046 4118
rect 9 3446 115076 4002
rect 9 3330 70 3446
rect 430 3330 115076 3446
rect 9 3110 115076 3330
rect 9 2994 115046 3110
rect 9 2102 115076 2994
rect 9 1986 70 2102
rect 430 1986 115076 2102
rect 9 1766 115076 1986
rect 9 1650 115046 1766
rect 9 1094 115076 1650
rect 9 978 70 1094
rect 430 978 115076 1094
rect 9 910 115076 978
<< metal4 >>
rect 2224 1538 2384 115670
rect 9904 1538 10064 115670
rect 17584 1538 17744 115670
rect 25264 1538 25424 115670
rect 32944 1538 33104 115670
rect 40624 1538 40784 115670
rect 48304 1538 48464 115670
rect 55984 1538 56144 115670
rect 63664 1538 63824 115670
rect 71344 1538 71504 115670
rect 79024 1538 79184 115670
rect 86704 1538 86864 115670
rect 94384 1538 94544 115670
rect 102064 1538 102224 115670
rect 109744 1538 109904 115670
<< obsm4 >>
rect 6174 1745 9874 115463
rect 10094 1745 17554 115463
rect 17774 1745 25234 115463
rect 25454 1745 32914 115463
rect 33134 1745 40594 115463
rect 40814 1745 48274 115463
rect 48494 1745 55954 115463
rect 56174 1745 63634 115463
rect 63854 1745 71314 115463
rect 71534 1745 78994 115463
rect 79214 1745 86674 115463
rect 86894 1745 94354 115463
rect 94574 1745 102034 115463
rect 102254 1745 109714 115463
rect 109934 1745 113946 115463
<< labels >>
rlabel metal2 s 67872 116868 67928 117168 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 14784 116868 14840 117168 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 88032 400 88088 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 115076 115920 115376 115976 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 7728 400 7784 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 85008 116868 85064 117168 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 115076 75264 115376 75320 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 100 54096 400 54152 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 115076 42336 115376 42392 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 100 116256 400 116312 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 113232 116868 113288 117168 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 100 92400 400 92456 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 115076 18816 115376 18872 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 100 59808 400 59864 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 24864 116868 24920 117168 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 100 103824 400 103880 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 99456 100 99512 400 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 115076 24528 115376 24584 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 112896 100 112952 400 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 5376 400 5432 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 114240 116868 114296 117168 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 58800 116868 58856 117168 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 100 12432 400 12488 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 100 22512 400 22568 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 55440 116868 55496 117168 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 115076 112560 115376 112616 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 12432 116868 12488 117168 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 115076 87696 115376 87752 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 100 66528 400 66584 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 98448 116868 98504 117168 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 115076 28896 115376 28952 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 100 40656 400 40712 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 115076 49392 115376 49448 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 9072 116868 9128 117168 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 94080 116868 94136 117168 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 40656 100 40712 400 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 115076 90048 115376 90104 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23520 100 23576 400 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 115076 10752 115376 10808 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 115076 19824 115376 19880 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 85680 100 85736 400 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 63504 116868 63560 117168 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 112896 400 112952 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 100 2016 400 2072 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 19488 116868 19544 117168 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 30576 116868 30632 117168 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 15792 116868 15848 117168 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 87024 400 87080 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 68880 100 68936 400 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 115076 101136 115376 101192 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 115076 25536 115376 25592 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 100 89040 400 89096 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 108192 100 108248 400 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 100 100464 400 100520 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 95760 100 95816 400 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 49728 116868 49784 117168 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 62160 116868 62216 117168 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 103824 100 103880 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 115076 41328 115376 41384 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 83664 116868 83720 117168 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 97440 116868 97496 117168 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 11088 100 11144 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 109872 116868 109928 117168 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 46032 100 46088 400 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 17136 116868 17192 117168 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 4704 116868 4760 117168 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 100 51744 400 51800 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 97104 100 97160 400 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 115076 46032 115376 46088 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 101808 116868 101864 117168 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 39312 400 39368 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 115076 17472 115376 17528 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 106512 116868 106568 117168 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 48384 100 48440 400 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 72240 100 72296 400 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 115076 13104 115376 13160 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 115076 72912 115376 72968 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 100 78960 400 79016 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 115076 105840 115376 105896 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 52080 116868 52136 117168 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 13440 100 13496 400 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 77952 400 78008 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 74592 100 74648 400 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 7728 100 7784 400 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 115076 66192 115376 66248 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 51744 100 51800 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 38304 100 38360 400 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 115076 37968 115376 38024 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98112 100 98168 400 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 108528 116868 108584 117168 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 115248 400 115304 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 100 60816 400 60872 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 76608 100 76664 400 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 65520 116868 65576 117168 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 100 73248 400 73304 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 115076 23184 115376 23240 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 100 44016 400 44072 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 100 53088 400 53144 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 75600 100 75656 400 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 115076 16464 115376 16520 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 115076 114912 115376 114968 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 115076 4032 115376 4088 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 26208 116868 26264 117168 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 56784 116868 56840 117168 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 100 48384 400 48440 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 67536 400 67592 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 71232 116868 71288 117168 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 83328 100 83384 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 10416 116868 10472 117168 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 34944 400 35000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 113904 100 113960 400 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 42672 100 42728 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 34944 100 35000 400 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 47712 116868 47768 117168 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 105168 116868 105224 117168 6 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 54096 100 54152 400 6 la_data_in[11]
port 117 nsew signal input
rlabel metal3 s 100 70896 400 70952 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 90384 116868 90440 117168 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 115076 113568 115376 113624 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 115076 29904 115376 29960 6 la_data_in[15]
port 121 nsew signal input
rlabel metal3 s 100 75600 400 75656 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 115076 22176 115376 22232 6 la_data_in[17]
port 123 nsew signal input
rlabel metal3 s 100 11088 400 11144 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 92736 116868 92792 117168 6 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 72576 116868 72632 117168 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 115076 96768 115376 96824 6 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 86016 116868 86072 117168 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 100 33600 400 33656 6 la_data_in[23]
port 130 nsew signal input
rlabel metal3 s 100 56448 400 56504 6 la_data_in[24]
port 131 nsew signal input
rlabel metal3 s 100 99456 400 99512 6 la_data_in[25]
port 132 nsew signal input
rlabel metal3 s 115076 106848 115376 106904 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 115076 63840 115376 63896 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 113904 400 113960 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 115076 48048 115376 48104 6 la_data_in[29]
port 136 nsew signal input
rlabel metal3 s 115076 100128 115376 100184 6 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 109536 100 109592 400 6 la_data_in[30]
port 138 nsew signal input
rlabel metal3 s 100 26880 400 26936 6 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 81312 100 81368 400 6 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 42000 116868 42056 117168 6 la_data_in[33]
port 141 nsew signal input
rlabel metal3 s 100 79968 400 80024 6 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 48720 116868 48776 117168 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 77952 116868 78008 117168 6 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 39312 100 39368 400 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 55104 100 55160 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal3 s 100 110544 400 110600 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 100 49728 400 49784 6 la_data_in[3]
port 148 nsew signal input
rlabel metal3 s 100 82320 400 82376 6 la_data_in[40]
port 149 nsew signal input
rlabel metal3 s 115076 84336 115376 84392 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 115076 83328 115376 83384 6 la_data_in[42]
port 151 nsew signal input
rlabel metal3 s 100 10080 400 10136 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 100 30240 400 30296 6 la_data_in[44]
port 153 nsew signal input
rlabel metal3 s 100 8736 400 8792 6 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 28224 100 28280 400 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 46368 116868 46424 117168 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 53088 100 53144 400 6 la_data_in[48]
port 157 nsew signal input
rlabel metal3 s 100 106176 400 106232 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 35280 116868 35336 117168 6 la_data_in[4]
port 159 nsew signal input
rlabel metal3 s 115076 31248 115376 31304 6 la_data_in[50]
port 160 nsew signal input
rlabel metal3 s 100 31584 400 31640 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 100 32592 400 32648 6 la_data_in[52]
port 162 nsew signal input
rlabel metal3 s 115076 3024 115376 3080 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 41664 100 41720 400 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 45024 400 45080 6 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 20160 100 20216 400 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 80304 116868 80360 117168 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 88368 116868 88424 117168 6 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 67536 100 67592 400 6 la_data_in[59]
port 169 nsew signal input
rlabel metal3 s 115076 56112 115376 56168 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 100 57456 400 57512 6 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 0 116868 56 117168 6 la_data_in[61]
port 172 nsew signal input
rlabel metal3 s 100 97104 400 97160 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 64512 116868 64568 117168 6 la_data_in[63]
port 174 nsew signal input
rlabel metal3 s 100 16800 400 16856 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 100 72240 400 72296 6 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 82320 100 82376 400 6 la_data_in[8]
port 177 nsew signal input
rlabel metal3 s 100 84672 400 84728 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 32928 116868 32984 117168 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 115076 47040 115376 47096 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 115076 109200 115376 109256 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 115076 62832 115376 62888 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 57792 116868 57848 117168 6 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 51072 116868 51128 117168 6 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 60816 100 60872 400 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 115076 53760 115376 53816 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 54432 116868 54488 117168 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 115076 80976 115376 81032 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 61152 116868 61208 117168 6 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 33600 100 33656 400 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 100 17808 400 17864 6 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 62160 100 62216 400 6 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 100800 116868 100856 117168 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 15792 100 15848 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 15792 400 15848 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 49728 100 49784 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 91392 400 91448 6 la_data_out[26]
port 197 nsew signal output
rlabel metal3 s 115076 52752 115376 52808 6 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 3360 116868 3416 117168 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 18144 116868 18200 117168 6 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 2352 116868 2408 117168 6 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 56448 100 56504 400 6 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 31584 100 31640 400 6 la_data_out[31]
port 203 nsew signal output
rlabel metal3 s 115076 93408 115376 93464 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 115076 44688 115376 44744 6 la_data_out[33]
port 205 nsew signal output
rlabel metal3 s 115076 1680 115376 1736 6 la_data_out[34]
port 206 nsew signal output
rlabel metal3 s 115076 15456 115376 15512 6 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 81648 116868 81704 117168 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 100 104832 400 104888 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 115076 34608 115376 34664 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 115076 97776 115376 97832 6 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 6720 100 6776 400 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 47376 100 47432 400 6 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 70224 116868 70280 117168 6 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 106176 100 106232 400 6 la_data_out[42]
port 215 nsew signal output
rlabel metal3 s 100 83328 400 83384 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 26880 100 26936 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 104832 100 104888 400 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 66864 116868 66920 117168 6 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 40656 116868 40712 117168 6 la_data_out[47]
port 220 nsew signal output
rlabel metal3 s 100 42672 400 42728 6 la_data_out[48]
port 221 nsew signal output
rlabel metal3 s 115076 7392 115376 7448 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 64176 100 64232 400 6 la_data_out[4]
port 223 nsew signal output
rlabel metal3 s 100 109536 400 109592 6 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 44352 116868 44408 117168 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 115076 26544 115376 26600 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 93744 400 93800 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 115076 79632 115376 79688 6 la_data_out[54]
port 228 nsew signal output
rlabel metal3 s 115076 103488 115376 103544 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 115076 69552 115376 69608 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 95088 116868 95144 117168 6 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 30240 100 30296 400 6 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 100464 100 100520 400 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 115076 8736 115376 8792 6 la_data_out[5]
port 234 nsew signal output
rlabel metal3 s 100 81312 400 81368 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 111888 116868 111944 117168 6 la_data_out[61]
port 236 nsew signal output
rlabel metal3 s 100 108192 400 108248 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 115076 54768 115376 54824 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 115076 43680 115376 43736 6 la_data_out[6]
port 239 nsew signal output
rlabel metal3 s 115076 81984 115376 82040 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 115076 65184 115376 65240 6 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 45360 116868 45416 117168 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 100 41664 400 41720 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 100 4368 400 4424 6 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 101472 100 101528 400 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 16800 100 16856 400 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 14448 400 14504 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 8064 116868 8120 117168 6 la_oenb[14]
port 248 nsew signal input
rlabel metal3 s 115076 9744 115376 9800 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 22848 116868 22904 117168 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 102816 400 102872 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 20496 116868 20552 117168 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 100 3360 400 3416 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 32592 100 32648 400 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 29232 400 29288 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 102816 100 102872 400 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 23856 116868 23912 117168 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 21168 100 21224 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 115076 60480 115376 60536 6 la_oenb[24]
port 259 nsew signal input
rlabel metal3 s 115076 110208 115376 110264 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 115248 116868 115304 117168 6 la_oenb[26]
port 261 nsew signal input
rlabel metal3 s 115076 99120 115376 99176 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 115076 95760 115376 95816 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 115076 94416 115376 94472 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 58464 100 58520 400 6 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 104160 116868 104216 117168 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 3360 100 3416 400 6 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 1008 100 1064 400 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 1344 116868 1400 117168 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 59808 100 59864 400 6 la_oenb[34]
port 270 nsew signal input
rlabel metal3 s 100 50736 400 50792 6 la_oenb[35]
port 271 nsew signal input
rlabel metal3 s 100 64176 400 64232 6 la_oenb[36]
port 272 nsew signal input
rlabel metal3 s 100 37296 400 37352 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 43008 116868 43064 117168 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 74592 400 74648 6 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 22512 100 22568 400 6 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 50736 100 50792 400 6 la_oenb[40]
port 277 nsew signal input
rlabel metal3 s 100 58464 400 58520 6 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 92400 100 92456 400 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 44016 100 44072 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal3 s 100 85680 400 85736 6 la_oenb[44]
port 281 nsew signal input
rlabel metal3 s 115076 57120 115376 57176 6 la_oenb[45]
port 282 nsew signal input
rlabel metal3 s 115076 77616 115376 77672 6 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 89040 100 89096 400 6 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 37296 116868 37352 117168 6 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 115248 100 115304 400 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 115076 74256 115376 74312 6 la_oenb[4]
port 287 nsew signal input
rlabel metal3 s 100 69888 400 69944 6 la_oenb[50]
port 288 nsew signal input
rlabel metal3 s 115076 59472 115376 59528 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 88032 100 88088 400 6 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 102816 116868 102872 117168 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 115076 12096 115376 12152 6 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 69216 116868 69272 117168 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 107184 100 107240 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 28224 116868 28280 117168 6 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 14448 100 14504 400 6 la_oenb[58]
port 296 nsew signal input
rlabel metal3 s 100 1008 400 1064 6 la_oenb[59]
port 297 nsew signal input
rlabel metal3 s 100 111888 400 111944 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 115076 76272 115376 76328 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 29232 100 29288 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 110544 100 110600 400 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 21168 400 21224 6 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 99456 116868 99512 117168 6 la_oenb[6]
port 303 nsew signal input
rlabel metal3 s 115076 88704 115376 88760 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 29568 116868 29624 117168 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 39648 116868 39704 117168 6 la_oenb[9]
port 306 nsew signal input
rlabel metal4 s 2224 1538 2384 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 115670 6 vdd
port 307 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 115670 6 vss
port 308 nsew ground bidirectional
rlabel metal3 s 115076 21168 115376 21224 6 wb_clk_i
port 309 nsew signal input
rlabel metal2 s 21504 116868 21560 117168 6 wb_rst_i
port 310 nsew signal input
rlabel metal3 s 115076 40320 115376 40376 6 wbs_ack_o
port 311 nsew signal output
rlabel metal2 s 76944 116868 77000 117168 6 wbs_adr_i[0]
port 312 nsew signal input
rlabel metal2 s 53088 116868 53144 117168 6 wbs_adr_i[10]
port 313 nsew signal input
rlabel metal2 s 7056 116868 7112 117168 6 wbs_adr_i[11]
port 314 nsew signal input
rlabel metal2 s 10080 100 10136 400 6 wbs_adr_i[12]
port 315 nsew signal input
rlabel metal3 s 100 28224 400 28280 6 wbs_adr_i[13]
port 316 nsew signal input
rlabel metal3 s 115076 85344 115376 85400 6 wbs_adr_i[14]
port 317 nsew signal input
rlabel metal3 s 115076 78624 115376 78680 6 wbs_adr_i[15]
port 318 nsew signal input
rlabel metal2 s 73248 100 73304 400 6 wbs_adr_i[16]
port 319 nsew signal input
rlabel metal3 s 100 65520 400 65576 6 wbs_adr_i[17]
port 320 nsew signal input
rlabel metal3 s 115076 36960 115376 37016 6 wbs_adr_i[18]
port 321 nsew signal input
rlabel metal2 s 111888 100 111944 400 6 wbs_adr_i[19]
port 322 nsew signal input
rlabel metal2 s 74592 116868 74648 117168 6 wbs_adr_i[1]
port 323 nsew signal input
rlabel metal3 s 100 63168 400 63224 6 wbs_adr_i[20]
port 324 nsew signal input
rlabel metal2 s 65520 100 65576 400 6 wbs_adr_i[21]
port 325 nsew signal input
rlabel metal2 s 93744 100 93800 400 6 wbs_adr_i[22]
port 326 nsew signal input
rlabel metal3 s 115076 27888 115376 27944 6 wbs_adr_i[23]
port 327 nsew signal input
rlabel metal2 s 13776 116868 13832 117168 6 wbs_adr_i[24]
port 328 nsew signal input
rlabel metal3 s 100 20160 400 20216 6 wbs_adr_i[25]
port 329 nsew signal input
rlabel metal2 s 12432 100 12488 400 6 wbs_adr_i[26]
port 330 nsew signal input
rlabel metal2 s 38640 116868 38696 117168 6 wbs_adr_i[27]
port 331 nsew signal input
rlabel metal3 s 115076 68544 115376 68600 6 wbs_adr_i[28]
port 332 nsew signal input
rlabel metal3 s 115076 111552 115376 111608 6 wbs_adr_i[29]
port 333 nsew signal input
rlabel metal3 s 100 13440 400 13496 6 wbs_adr_i[2]
port 334 nsew signal input
rlabel metal3 s 100 46032 400 46088 6 wbs_adr_i[30]
port 335 nsew signal input
rlabel metal3 s 115076 50400 115376 50456 6 wbs_adr_i[31]
port 336 nsew signal input
rlabel metal2 s 90384 100 90440 400 6 wbs_adr_i[3]
port 337 nsew signal input
rlabel metal2 s 89376 116868 89432 117168 6 wbs_adr_i[4]
port 338 nsew signal input
rlabel metal2 s 87024 100 87080 400 6 wbs_adr_i[5]
port 339 nsew signal input
rlabel metal2 s 37296 100 37352 400 6 wbs_adr_i[6]
port 340 nsew signal input
rlabel metal2 s 5376 100 5432 400 6 wbs_adr_i[7]
port 341 nsew signal input
rlabel metal3 s 115076 672 115376 728 6 wbs_adr_i[8]
port 342 nsew signal input
rlabel metal3 s 115076 32256 115376 32312 6 wbs_adr_i[9]
port 343 nsew signal input
rlabel metal2 s 36288 116868 36344 117168 6 wbs_cyc_i
port 344 nsew signal input
rlabel metal3 s 115076 102480 115376 102536 6 wbs_dat_i[0]
port 345 nsew signal input
rlabel metal3 s 100 90384 400 90440 6 wbs_dat_i[10]
port 346 nsew signal input
rlabel metal3 s 100 98112 400 98168 6 wbs_dat_i[11]
port 347 nsew signal input
rlabel metal3 s 100 94752 400 94808 6 wbs_dat_i[12]
port 348 nsew signal input
rlabel metal2 s 4368 100 4424 400 6 wbs_dat_i[13]
port 349 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 wbs_dat_i[14]
port 350 nsew signal input
rlabel metal3 s 115076 61824 115376 61880 6 wbs_dat_i[15]
port 351 nsew signal input
rlabel metal2 s 66528 100 66584 400 6 wbs_dat_i[16]
port 352 nsew signal input
rlabel metal3 s 100 19152 400 19208 6 wbs_dat_i[17]
port 353 nsew signal input
rlabel metal2 s 107520 116868 107576 117168 6 wbs_dat_i[18]
port 354 nsew signal input
rlabel metal2 s 5712 116868 5768 117168 6 wbs_dat_i[19]
port 355 nsew signal input
rlabel metal2 s 17808 100 17864 400 6 wbs_dat_i[1]
port 356 nsew signal input
rlabel metal3 s 115076 70896 115376 70952 6 wbs_dat_i[20]
port 357 nsew signal input
rlabel metal2 s 110880 116868 110936 117168 6 wbs_dat_i[21]
port 358 nsew signal input
rlabel metal3 s 100 68880 400 68936 6 wbs_dat_i[22]
port 359 nsew signal input
rlabel metal3 s 115076 92064 115376 92120 6 wbs_dat_i[23]
port 360 nsew signal input
rlabel metal3 s 115076 38976 115376 39032 6 wbs_dat_i[24]
port 361 nsew signal input
rlabel metal2 s 79968 100 80024 400 6 wbs_dat_i[25]
port 362 nsew signal input
rlabel metal2 s 96096 116868 96152 117168 6 wbs_dat_i[26]
port 363 nsew signal input
rlabel metal2 s 27216 116868 27272 117168 6 wbs_dat_i[27]
port 364 nsew signal input
rlabel metal2 s 35952 100 36008 400 6 wbs_dat_i[28]
port 365 nsew signal input
rlabel metal3 s 115076 71904 115376 71960 6 wbs_dat_i[29]
port 366 nsew signal input
rlabel metal2 s 94752 100 94808 400 6 wbs_dat_i[2]
port 367 nsew signal input
rlabel metal3 s 115076 35616 115376 35672 6 wbs_dat_i[30]
port 368 nsew signal input
rlabel metal3 s 100 62160 400 62216 6 wbs_dat_i[31]
port 369 nsew signal input
rlabel metal3 s 115076 5040 115376 5096 6 wbs_dat_i[3]
port 370 nsew signal input
rlabel metal2 s 19152 100 19208 400 6 wbs_dat_i[4]
port 371 nsew signal input
rlabel metal2 s 57456 100 57512 400 6 wbs_dat_i[5]
port 372 nsew signal input
rlabel metal3 s 115076 51408 115376 51464 6 wbs_dat_i[6]
port 373 nsew signal input
rlabel metal2 s 91728 116868 91784 117168 6 wbs_dat_i[7]
port 374 nsew signal input
rlabel metal3 s 115076 104496 115376 104552 6 wbs_dat_i[8]
port 375 nsew signal input
rlabel metal3 s 115076 6384 115376 6440 6 wbs_dat_i[9]
port 376 nsew signal input
rlabel metal3 s 100 23520 400 23576 6 wbs_dat_o[0]
port 377 nsew signal output
rlabel metal3 s 115076 67200 115376 67256 6 wbs_dat_o[10]
port 378 nsew signal output
rlabel metal2 s 2016 100 2072 400 6 wbs_dat_o[11]
port 379 nsew signal output
rlabel metal3 s 115076 108192 115376 108248 6 wbs_dat_o[12]
port 380 nsew signal output
rlabel metal2 s 87024 116868 87080 117168 6 wbs_dat_o[13]
port 381 nsew signal output
rlabel metal3 s 115076 14112 115376 14168 6 wbs_dat_o[14]
port 382 nsew signal output
rlabel metal2 s 82656 116868 82712 117168 6 wbs_dat_o[15]
port 383 nsew signal output
rlabel metal2 s 78960 100 79016 400 6 wbs_dat_o[16]
port 384 nsew signal output
rlabel metal3 s 100 35952 400 36008 6 wbs_dat_o[17]
port 385 nsew signal output
rlabel metal2 s 77952 100 78008 400 6 wbs_dat_o[18]
port 386 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 387 nsew signal output
rlabel metal2 s 91392 100 91448 400 6 wbs_dat_o[1]
port 388 nsew signal output
rlabel metal3 s 100 55104 400 55160 6 wbs_dat_o[20]
port 389 nsew signal output
rlabel metal3 s 100 101472 400 101528 6 wbs_dat_o[21]
port 390 nsew signal output
rlabel metal2 s 31920 116868 31976 117168 6 wbs_dat_o[22]
port 391 nsew signal output
rlabel metal3 s 100 38304 400 38360 6 wbs_dat_o[23]
port 392 nsew signal output
rlabel metal2 s 24864 100 24920 400 6 wbs_dat_o[24]
port 393 nsew signal output
rlabel metal2 s 8736 100 8792 400 6 wbs_dat_o[25]
port 394 nsew signal output
rlabel metal2 s 60144 116868 60200 117168 6 wbs_dat_o[26]
port 395 nsew signal output
rlabel metal2 s 33936 116868 33992 117168 6 wbs_dat_o[27]
port 396 nsew signal output
rlabel metal2 s 63168 100 63224 400 6 wbs_dat_o[28]
port 397 nsew signal output
rlabel metal2 s 79296 116868 79352 117168 6 wbs_dat_o[29]
port 398 nsew signal output
rlabel metal3 s 115076 33600 115376 33656 6 wbs_dat_o[2]
port 399 nsew signal output
rlabel metal3 s 100 76608 400 76664 6 wbs_dat_o[30]
port 400 nsew signal output
rlabel metal3 s 115076 91056 115376 91112 6 wbs_dat_o[31]
port 401 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 wbs_dat_o[3]
port 402 nsew signal output
rlabel metal2 s 45024 100 45080 400 6 wbs_dat_o[4]
port 403 nsew signal output
rlabel metal2 s 69888 100 69944 400 6 wbs_dat_o[5]
port 404 nsew signal output
rlabel metal3 s 115076 86688 115376 86744 6 wbs_dat_o[6]
port 405 nsew signal output
rlabel metal2 s 70896 100 70952 400 6 wbs_dat_o[7]
port 406 nsew signal output
rlabel metal2 s 75936 116868 75992 117168 6 wbs_dat_o[8]
port 407 nsew signal output
rlabel metal2 s 73584 116868 73640 117168 6 wbs_dat_o[9]
port 408 nsew signal output
rlabel metal3 s 100 107184 400 107240 6 wbs_sel_i[0]
port 409 nsew signal input
rlabel metal2 s 11424 116868 11480 117168 6 wbs_sel_i[1]
port 410 nsew signal input
rlabel metal2 s 84672 100 84728 400 6 wbs_sel_i[2]
port 411 nsew signal input
rlabel metal3 s 100 25872 400 25928 6 wbs_sel_i[3]
port 412 nsew signal input
rlabel metal3 s 100 95760 400 95816 6 wbs_stb_i
port 413 nsew signal input
rlabel metal3 s 115076 58464 115376 58520 6 wbs_we_i
port 414 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 115476 117268
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35544274
string GDS_FILE /home/vijayan/CARAVEL_FLOW/GFmpw0/AES128_GFMPW0/openlane/aes_core/runs/22_11_28_10_11/results/signoff/aes_core.magic.gds
string GDS_START 457756
<< end >>

